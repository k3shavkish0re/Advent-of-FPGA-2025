`timescale 1ns/1ns

module tb_puzzle1;

    localparam int NUM_BANKS = 200;
    localparam int SIZE_BANK = 128;
    localparam int EFFECTIVE_DEPTH = 100;

    logic clk;
    logic rst_n;
    logic bank_en;
    logic [NUM_BANKS-1:0][3:0] val;
    logic [14:0] max_joltage;

    // Instantiate DUT
    puzzle1 #(
        .NUM_BANKS(NUM_BANKS),
        .SIZE_BANK(SIZE_BANK)
    ) dut (
        .clk(clk),
        .rst_n(rst_n),
        .bank_en(bank_en),
        .val(val),
        .max_joltage(max_joltage)
    );
	
	// ----------------------------------------
    // $monitor — print internal DUT signals
    // ----------------------------------------
    initial begin
        $monitor("[%0t] clk=%0b | rst_n=%0b | bank_en=%0d |state=%0d | bank_idx=%0d | cnt=%0d | sum=%0d | max_joltage=%0d",
            $time,
			clk,
			rst_n,
			bank_en,
            dut.state_q,
            dut.bank_index_cnt_q,
            dut.cnt_q,
            dut.sum_q,
            dut.max_joltage
        );
    end
	
	
	    final begin
            // Print all 200 banks
            for (int i = 0; i < 200; i++) begin
                $display("Bank[%0d]: max=%0d",
                        i,
                        dut.max_in_bank_q[i]
                );
            end
            $display("---------------------------------------------------------");
        end
	
	
	
	
    // Clock
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    initial begin
        $dumpfile("tb.vcd");
        $dumpvars(0, tb_puzzle1);

        rst_n  = 1;
        bank_en = 0;
        val     = '0;

        repeat (5) @(posedge clk);
        rst_n = 0;
        repeat (5) @(posedge clk);
        rst_n = 1;
        @(posedge clk);

        // Start storing
        bank_en = 1;
        @(posedge clk);
        bank_en = 1;   // keep high during storage

        // ---------------- INPUT-DRIVEN VAL PATTERN ----------------
        val = '{ 7, 5, 2, 4, 1, 5, 3, 2, 5, 4, 5, 6, 2, 2, 4, 6, 1, 4, 5, 9, 2, 2, 3, 2, 3, 4, 1, 3, 6, 2, 3, 4, 1, 3, 1, 4, 2, 3, 8, 4, 2, 5, 5, 2, 5, 4, 6, 1, 3, 2, 1, 2, 4, 2, 1, 1, 3, 2, 2, 5, 7, 1, 5, 7, 3, 5, 3, 5, 2, 3, 2, 3, 5, 4, 1, 3, 4, 2, 2, 1, 3, 3, 4, 9, 2, 3, 1, 4, 3, 4, 3, 4, 2, 4, 2, 3, 3, 5, 4, 1, 3, 5, 2, 1, 3, 3, 6, 2, 2, 3, 4, 3, 4, 2, 4, 3, 6, 3, 6, 2, 4, 4, 1, 1, 4, 2, 3, 8, 7, 4, 4, 2, 4, 6, 3, 3, 4, 7, 5, 2, 3, 3, 3, 3, 2, 2, 2, 2, 2, 1, 7, 2, 3, 2, 7, 3, 2, 4, 6, 2, 3, 3, 3, 2, 7, 4, 3, 5, 1, 3, 4, 5, 3, 7, 5, 8, 2, 4, 3, 3, 5, 1, 5, 3, 6, 2, 2, 3, 3, 1, 4, 3, 1, 3, 2, 5, 2, 5, 2, 2 };
        @(posedge clk);
        val = '{ 3, 4, 3, 3, 2, 4, 2, 3, 6, 2, 4, 5, 3, 2, 1, 3, 3, 2, 3, 2, 2, 2, 5, 2, 3, 2, 1, 7, 6, 2, 3, 4, 2, 3, 4, 5, 1, 2, 2, 5, 2, 4, 8, 7, 4, 4, 4, 1, 1, 2, 6, 1, 4, 2, 2, 2, 2, 2, 4, 4, 3, 4, 4, 9, 3, 2, 6, 4, 2, 4, 1, 3, 1, 9, 3, 2, 4, 1, 5, 3, 3, 2, 2, 6, 2, 6, 2, 2, 3, 2, 5, 4, 4, 2, 5, 3, 7, 1, 5, 3, 7, 5, 3, 7, 4, 6, 4, 4, 3, 6, 2, 3, 2, 4, 2, 2, 2, 5, 2, 2, 4, 3, 3, 2, 2, 5, 1, 6, 5, 4, 7, 2, 2, 2, 4, 2, 2, 4, 3, 2, 1, 3, 3, 1, 4, 3, 2, 2, 2, 2, 4, 3, 4, 2, 4, 3, 6, 1, 2, 2, 4, 2, 2, 2, 3, 5, 5, 4, 5, 9, 4, 3, 5, 4, 3, 8, 9, 4, 4, 1, 4, 2, 8, 2, 2, 2, 2, 2, 2, 2, 6, 4, 3, 2, 2, 7, 2, 3, 1, 2 };
        @(posedge clk);
        val = '{ 5, 3, 4, 3, 3, 7, 7, 1, 4, 4, 4, 4, 2, 3, 4, 5, 2, 1, 5, 2, 3, 1, 4, 2, 2, 2, 2, 5, 6, 2, 2, 2, 2, 2, 3, 4, 2, 3, 2, 6, 1, 5, 4, 9, 5, 4, 3, 3, 5, 2, 4, 4, 4, 2, 3, 3, 2, 2, 2, 3, 5, 3, 1, 4, 1, 2, 8, 9, 4, 3, 2, 3, 2, 5, 5, 4, 3, 2, 3, 3, 2, 3, 2, 6, 3, 9, 1, 3, 3, 4, 8, 3, 1, 3, 3, 5, 3, 6, 2, 3, 2, 5, 4, 2, 5, 5, 5, 4, 5, 5, 2, 3, 4, 2, 3, 2, 2, 6, 7, 4, 2, 3, 2, 2, 3, 2, 6, 8, 3, 6, 8, 4, 2, 8, 1, 3, 3, 4, 4, 6, 2, 3, 8, 3, 6, 4, 2, 3, 3, 2, 4, 4, 3, 5, 1, 5, 4, 3, 2, 2, 2, 2, 2, 2, 6, 2, 5, 4, 4, 2, 2, 3, 5, 4, 5, 7, 1, 7, 1, 2, 2, 1, 2, 3, 7, 1, 2, 9, 7, 4, 7, 4, 2, 1, 2, 4, 3, 1, 1, 2 };
        @(posedge clk);
        val = '{ 1, 3, 4, 1, 3, 5, 6, 2, 7, 4, 3, 4, 2, 2, 2, 3, 3, 1, 4, 2, 1, 3, 4, 3, 3, 2, 4, 4, 7, 2, 2, 3, 4, 3, 2, 8, 2, 1, 8, 4, 1, 6, 2, 5, 2, 2, 3, 1, 2, 2, 2, 1, 4, 4, 7, 1, 3, 2, 2, 4, 2, 2, 5, 7, 3, 1, 5, 5, 6, 4, 6, 4, 4, 5, 4, 9, 3, 1, 2, 2, 3, 5, 2, 7, 2, 1, 1, 8, 3, 5, 3, 6, 4, 3, 2, 5, 7, 5, 2, 2, 4, 7, 3, 2, 2, 4, 6, 1, 4, 6, 3, 3, 1, 2, 4, 4, 2, 6, 3, 1, 2, 2, 6, 2, 4, 3, 6, 9, 9, 4, 1, 4, 3, 6, 3, 1, 2, 5, 2, 9, 2, 3, 2, 2, 2, 2, 3, 3, 3, 2, 2, 4, 3, 4, 6, 4, 2, 4, 2, 8, 2, 3, 4, 2, 7, 3, 4, 3, 2, 1, 3, 2, 3, 6, 4, 5, 2, 1, 2, 3, 2, 2, 2, 2, 3, 2, 4, 4, 3, 4, 4, 1, 1, 2, 2, 5, 4, 1, 3, 2 };
        @(posedge clk);
        val = '{ 2, 4, 3, 2, 3, 4, 3, 2, 5, 4, 4, 4, 2, 1, 2, 2, 4, 4, 4, 2, 3, 3, 3, 1, 2, 8, 5, 1, 3, 2, 2, 4, 4, 2, 3, 5, 3, 3, 3, 5, 3, 5, 5, 7, 2, 4, 4, 5, 5, 2, 6, 2, 6, 4, 8, 2, 2, 2, 3, 3, 4, 3, 2, 5, 5, 2, 3, 2, 5, 4, 6, 1, 2, 7, 4, 9, 3, 3, 4, 3, 4, 2, 2, 5, 5, 4, 2, 3, 3, 4, 5, 7, 3, 3, 1, 5, 3, 4, 1, 2, 1, 2, 2, 5, 5, 4, 3, 2, 4, 4, 2, 3, 1, 2, 3, 2, 3, 1, 5, 5, 3, 2, 2, 2, 2, 4, 5, 4, 7, 2, 7, 6, 3, 2, 4, 3, 2, 4, 2, 1, 5, 3, 1, 1, 2, 1, 2, 5, 3, 1, 3, 4, 3, 2, 8, 3, 7, 5, 2, 3, 1, 2, 2, 1, 7, 3, 3, 5, 2, 4, 3, 2, 1, 6, 5, 5, 2, 3, 4, 4, 3, 3, 1, 3, 3, 2, 2, 3, 2, 4, 5, 2, 2, 2, 2, 1, 3, 4, 3, 4 };
        @(posedge clk);
        val = '{ 3, 4, 2, 3, 2, 4, 2, 2, 6, 4, 4, 5, 2, 1, 2, 1, 5, 4, 4, 1, 2, 4, 8, 1, 2, 2, 6, 3, 7, 2, 2, 3, 2, 4, 3, 4, 6, 8, 5, 4, 2, 6, 2, 7, 3, 2, 3, 5, 5, 2, 3, 2, 9, 2, 2, 1, 3, 2, 3, 4, 6, 4, 2, 9, 2, 2, 4, 7, 5, 5, 2, 4, 2, 4, 2, 2, 3, 2, 4, 3, 3, 4, 2, 5, 2, 2, 6, 5, 3, 2, 3, 2, 4, 1, 6, 6, 2, 5, 5, 2, 5, 3, 3, 4, 6, 3, 6, 6, 1, 4, 2, 4, 2, 2, 3, 2, 4, 3, 4, 2, 3, 3, 4, 1, 4, 1, 6, 6, 8, 5, 5, 2, 1, 6, 2, 2, 2, 4, 1, 2, 3, 2, 2, 3, 1, 2, 2, 1, 3, 1, 4, 2, 2, 4, 2, 4, 2, 5, 2, 2, 3, 1, 4, 2, 5, 1, 4, 6, 3, 6, 4, 4, 4, 7, 3, 7, 2, 3, 2, 2, 2, 6, 2, 3, 3, 2, 1, 8, 3, 2, 5, 2, 2, 2, 3, 2, 4, 7, 2, 1 };
        @(posedge clk);
        val = '{ 3, 5, 3, 3, 3, 3, 2, 2, 6, 4, 6, 5, 2, 1, 4, 6, 3, 1, 8, 4, 4, 4, 2, 2, 3, 4, 1, 6, 6, 4, 2, 3, 1, 3, 6, 7, 1, 2, 2, 8, 2, 6, 6, 5, 5, 7, 4, 4, 7, 3, 5, 3, 4, 4, 4, 1, 2, 2, 2, 4, 9, 4, 3, 5, 1, 3, 7, 3, 2, 2, 5, 4, 2, 5, 5, 5, 4, 2, 4, 3, 3, 2, 2, 9, 2, 4, 4, 2, 2, 2, 3, 8, 4, 1, 4, 1, 2, 5, 3, 2, 4, 1, 8, 5, 3, 4, 8, 3, 5, 7, 3, 3, 5, 2, 3, 2, 4, 5, 4, 2, 4, 2, 2, 2, 5, 1, 6, 4, 5, 7, 3, 2, 6, 3, 3, 3, 2, 4, 1, 5, 3, 3, 1, 2, 3, 2, 1, 2, 6, 2, 3, 3, 5, 4, 8, 2, 3, 1, 5, 3, 3, 5, 3, 2, 6, 3, 9, 2, 1, 3, 7, 2, 3, 7, 2, 6, 2, 3, 2, 2, 6, 3, 3, 4, 2, 2, 2, 5, 5, 3, 6, 4, 2, 2, 1, 7, 5, 4, 1, 4 };
        @(posedge clk);
        val = '{ 2, 5, 2, 2, 2, 7, 3, 3, 9, 4, 5, 2, 2, 2, 8, 3, 3, 4, 5, 1, 3, 2, 3, 2, 3, 1, 3, 5, 4, 2, 2, 3, 1, 1, 3, 5, 7, 2, 4, 5, 2, 4, 4, 7, 5, 2, 4, 4, 2, 2, 3, 3, 4, 4, 6, 2, 2, 2, 5, 5, 4, 4, 3, 5, 3, 1, 6, 5, 2, 7, 5, 3, 2, 6, 4, 8, 2, 2, 1, 2, 4, 1, 4, 6, 6, 4, 1, 4, 2, 2, 2, 7, 2, 3, 2, 3, 2, 4, 3, 3, 6, 8, 7, 4, 3, 3, 3, 4, 3, 6, 4, 2, 3, 3, 3, 3, 4, 7, 3, 7, 3, 2, 3, 2, 9, 1, 6, 6, 8, 4, 7, 4, 2, 3, 3, 4, 4, 5, 3, 2, 5, 1, 2, 3, 4, 1, 3, 2, 2, 2, 3, 5, 4, 2, 6, 7, 2, 6, 4, 5, 2, 6, 2, 3, 4, 4, 2, 7, 2, 4, 2, 4, 4, 4, 5, 9, 1, 2, 4, 4, 6, 5, 4, 3, 6, 2, 2, 3, 3, 3, 4, 2, 1, 4, 2, 2, 2, 3, 6, 4 };
        @(posedge clk);
        val = '{ 3, 2, 5, 4, 2, 5, 3, 1, 4, 1, 5, 3, 2, 4, 2, 4, 4, 2, 9, 2, 2, 3, 2, 3, 5, 3, 2, 4, 3, 2, 2, 4, 1, 3, 3, 3, 4, 2, 5, 5, 3, 4, 4, 2, 4, 4, 3, 4, 5, 1, 6, 3, 5, 8, 5, 2, 1, 2, 2, 3, 5, 7, 4, 5, 4, 1, 6, 2, 1, 3, 6, 1, 2, 6, 3, 3, 2, 2, 3, 4, 3, 2, 2, 7, 2, 3, 3, 3, 7, 4, 2, 6, 4, 5, 2, 8, 2, 3, 2, 3, 6, 1, 3, 6, 3, 3, 3, 3, 3, 7, 2, 3, 2, 2, 3, 3, 5, 6, 6, 2, 5, 3, 4, 2, 7, 2, 7, 6, 5, 3, 3, 5, 2, 3, 4, 4, 4, 5, 4, 2, 3, 3, 2, 2, 2, 2, 1, 2, 8, 4, 4, 3, 4, 2, 3, 6, 3, 6, 3, 2, 3, 2, 4, 4, 4, 2, 4, 5, 2, 3, 4, 3, 4, 3, 5, 7, 2, 3, 3, 2, 4, 2, 5, 3, 3, 2, 2, 7, 2, 3, 5, 6, 2, 2, 2, 4, 5, 5, 2, 4 };
        @(posedge clk);
        val = '{ 2, 5, 4, 3, 3, 4, 3, 2, 2, 2, 4, 6, 1, 2, 6, 4, 2, 2, 4, 2, 5, 2, 5, 1, 5, 4, 7, 5, 4, 2, 1, 3, 4, 2, 2, 9, 5, 2, 2, 6, 1, 4, 7, 3, 2, 4, 5, 6, 3, 3, 2, 2, 3, 3, 6, 1, 1, 3, 3, 5, 2, 4, 1, 7, 5, 2, 3, 7, 6, 7, 7, 4, 3, 9, 3, 7, 3, 2, 4, 7, 1, 5, 2, 6, 5, 2, 7, 5, 2, 2, 1, 4, 4, 2, 7, 9, 2, 5, 2, 2, 1, 3, 3, 1, 3, 5, 6, 4, 4, 6, 3, 3, 4, 2, 3, 2, 2, 8, 3, 3, 4, 5, 9, 2, 6, 2, 6, 4, 7, 1, 5, 5, 5, 5, 3, 3, 2, 5, 3, 4, 9, 3, 2, 2, 2, 2, 2, 3, 3, 3, 5, 1, 2, 3, 7, 7, 3, 6, 2, 3, 1, 2, 2, 1, 4, 3, 3, 7, 2, 2, 7, 1, 6, 1, 7, 6, 2, 3, 1, 2, 3, 8, 1, 3, 4, 1, 1, 4, 3, 3, 3, 5, 3, 2, 1, 6, 4, 3, 2, 1 };
        @(posedge clk);
        val = '{ 2, 4, 2, 2, 3, 4, 3, 4, 4, 1, 3, 3, 1, 2, 1, 3, 3, 5, 4, 7, 5, 5, 4, 1, 2, 2, 3, 8, 6, 1, 2, 2, 3, 2, 2, 2, 3, 2, 1, 5, 1, 6, 3, 6, 4, 4, 3, 2, 3, 2, 6, 2, 4, 4, 3, 2, 2, 1, 2, 3, 7, 2, 1, 4, 2, 2, 4, 5, 5, 3, 3, 2, 2, 5, 2, 3, 5, 1, 4, 1, 4, 4, 2, 8, 5, 3, 1, 4, 3, 3, 8, 7, 2, 3, 2, 3, 1, 4, 2, 3, 3, 5, 1, 5, 3, 2, 4, 4, 3, 6, 3, 3, 2, 2, 3, 5, 3, 2, 2, 6, 4, 3, 5, 3, 7, 2, 5, 8, 8, 3, 3, 2, 4, 5, 3, 3, 2, 3, 2, 1, 3, 3, 2, 2, 5, 1, 3, 8, 9, 1, 5, 4, 2, 5, 3, 2, 2, 2, 2, 7, 5, 2, 2, 3, 6, 4, 3, 6, 2, 4, 4, 2, 5, 5, 5, 4, 2, 4, 2, 2, 5, 2, 2, 6, 7, 2, 3, 6, 3, 3, 6, 2, 2, 2, 5, 6, 5, 3, 3, 2 };
        @(posedge clk);
        val = '{ 2, 4, 3, 3, 3, 6, 3, 8, 7, 4, 4, 5, 2, 5, 7, 3, 4, 2, 5, 2, 2, 5, 4, 4, 2, 3, 2, 2, 4, 2, 2, 3, 3, 2, 2, 3, 1, 6, 3, 6, 2, 5, 3, 6, 5, 2, 3, 3, 7, 2, 3, 8, 3, 5, 2, 2, 2, 1, 2, 4, 4, 3, 4, 8, 1, 2, 4, 4, 3, 3, 6, 1, 2, 3, 4, 2, 3, 2, 3, 3, 5, 2, 4, 6, 3, 4, 3, 5, 4, 3, 4, 3, 4, 2, 2, 3, 6, 5, 2, 3, 3, 6, 1, 5, 3, 5, 6, 3, 2, 8, 3, 2, 3, 3, 3, 2, 7, 6, 6, 3, 4, 2, 2, 1, 4, 2, 5, 4, 4, 6, 4, 2, 2, 3, 3, 2, 3, 5, 2, 2, 2, 3, 1, 3, 8, 2, 1, 2, 3, 2, 4, 1, 6, 3, 4, 5, 1, 4, 2, 2, 1, 1, 3, 2, 5, 3, 1, 6, 2, 3, 7, 3, 4, 6, 3, 2, 3, 5, 1, 2, 4, 2, 2, 7, 7, 2, 2, 4, 1, 2, 6, 1, 2, 2, 1, 5, 4, 4, 5, 2 };
        @(posedge clk);
        val = '{ 3, 3, 8, 4, 3, 3, 2, 1, 8, 1, 6, 6, 4, 2, 2, 3, 3, 4, 4, 1, 3, 3, 4, 2, 4, 2, 7, 5, 4, 5, 3, 1, 3, 2, 2, 3, 1, 2, 4, 4, 2, 6, 5, 2, 2, 2, 2, 3, 2, 2, 3, 3, 6, 6, 2, 2, 3, 2, 2, 2, 2, 2, 3, 4, 3, 1, 9, 7, 2, 3, 6, 3, 3, 5, 5, 3, 3, 2, 3, 2, 1, 3, 2, 5, 5, 4, 3, 3, 3, 4, 8, 5, 5, 9, 4, 6, 3, 5, 1, 3, 5, 5, 2, 5, 2, 3, 6, 2, 4, 7, 3, 3, 1, 2, 4, 4, 2, 1, 3, 5, 2, 2, 4, 9, 4, 3, 4, 4, 9, 5, 4, 4, 1, 4, 3, 5, 1, 7, 1, 2, 5, 6, 1, 4, 4, 1, 2, 2, 3, 3, 4, 5, 4, 3, 5, 9, 2, 5, 5, 2, 3, 3, 3, 2, 3, 4, 2, 4, 2, 4, 3, 2, 3, 4, 6, 8, 2, 4, 2, 2, 2, 2, 1, 4, 2, 2, 3, 4, 2, 2, 5, 2, 2, 2, 2, 6, 3, 5, 3, 4 };
        @(posedge clk);
        val = '{ 3, 5, 3, 1, 2, 4, 3, 2, 4, 4, 6, 4, 1, 3, 7, 4, 2, 2, 7, 4, 2, 2, 4, 2, 2, 2, 8, 7, 5, 3, 1, 3, 3, 4, 2, 2, 4, 1, 6, 5, 2, 6, 5, 5, 4, 5, 6, 4, 2, 3, 2, 2, 3, 2, 2, 3, 7, 2, 7, 2, 2, 4, 1, 6, 3, 3, 3, 5, 6, 1, 6, 4, 2, 5, 8, 3, 4, 2, 4, 2, 3, 4, 1, 9, 2, 2, 6, 3, 1, 3, 2, 3, 4, 1, 5, 3, 2, 4, 3, 2, 8, 2, 2, 4, 5, 4, 7, 2, 2, 7, 4, 3, 2, 2, 4, 2, 5, 7, 5, 2, 3, 2, 4, 2, 6, 2, 5, 5, 8, 1, 3, 2, 5, 3, 3, 3, 2, 4, 4, 6, 6, 3, 2, 4, 1, 2, 2, 2, 3, 2, 3, 3, 1, 2, 1, 6, 3, 4, 2, 3, 2, 1, 5, 2, 5, 3, 3, 3, 3, 3, 6, 4, 3, 3, 4, 4, 3, 3, 2, 2, 2, 2, 5, 5, 2, 2, 1, 6, 5, 2, 3, 3, 1, 2, 2, 3, 4, 3, 2, 3 };
        @(posedge clk);
        val = '{ 2, 4, 2, 2, 5, 5, 5, 5, 3, 3, 6, 6, 2, 2, 3, 6, 3, 2, 5, 2, 2, 5, 3, 2, 2, 3, 1, 8, 2, 4, 3, 4, 2, 1, 3, 3, 3, 4, 2, 2, 3, 8, 5, 7, 2, 9, 6, 3, 3, 2, 4, 2, 4, 2, 6, 2, 3, 4, 2, 1, 2, 2, 3, 6, 3, 2, 3, 5, 3, 3, 4, 3, 4, 5, 1, 3, 1, 2, 1, 1, 6, 2, 2, 4, 7, 5, 2, 4, 2, 3, 6, 7, 4, 3, 5, 3, 6, 5, 3, 1, 5, 7, 3, 2, 3, 2, 5, 2, 2, 7, 7, 3, 3, 2, 2, 4, 6, 5, 5, 3, 4, 2, 2, 2, 4, 2, 4, 7, 8, 5, 6, 2, 1, 4, 4, 3, 2, 4, 2, 2, 2, 3, 2, 6, 9, 2, 2, 1, 3, 4, 4, 2, 3, 2, 2, 9, 3, 1, 2, 8, 3, 2, 3, 1, 7, 3, 3, 7, 3, 5, 2, 1, 4, 4, 4, 6, 2, 2, 5, 5, 4, 2, 2, 3, 1, 2, 2, 2, 3, 3, 3, 2, 3, 2, 2, 5, 7, 3, 6, 4 };
        @(posedge clk);
        val = '{ 2, 4, 4, 4, 3, 6, 3, 2, 6, 3, 4, 1, 2, 2, 7, 3, 4, 1, 7, 2, 3, 5, 9, 2, 3, 2, 2, 4, 7, 2, 2, 2, 2, 2, 2, 5, 6, 4, 3, 9, 5, 4, 6, 4, 4, 3, 2, 5, 2, 2, 3, 2, 2, 3, 6, 3, 2, 1, 2, 6, 3, 4, 3, 4, 3, 3, 4, 5, 4, 9, 7, 1, 2, 6, 5, 6, 4, 2, 2, 3, 1, 4, 1, 5, 6, 2, 1, 4, 1, 3, 5, 6, 3, 1, 3, 3, 6, 3, 2, 2, 3, 5, 2, 4, 3, 3, 8, 2, 3, 3, 4, 4, 2, 3, 3, 4, 5, 6, 6, 3, 2, 2, 9, 2, 2, 3, 5, 9, 4, 4, 6, 6, 2, 4, 5, 3, 1, 5, 3, 2, 1, 3, 2, 3, 4, 2, 2, 2, 6, 1, 4, 3, 3, 2, 8, 4, 4, 4, 4, 5, 3, 2, 2, 2, 6, 1, 5, 5, 2, 3, 6, 2, 3, 5, 3, 7, 4, 4, 2, 2, 5, 1, 1, 3, 6, 2, 1, 4, 3, 3, 4, 1, 2, 2, 3, 4, 2, 7, 6, 5 };
        @(posedge clk);
        val = '{ 5, 9, 3, 3, 2, 4, 3, 2, 8, 3, 6, 3, 2, 5, 6, 3, 2, 2, 3, 2, 3, 2, 4, 2, 4, 2, 3, 2, 4, 2, 3, 4, 1, 2, 2, 2, 3, 4, 3, 5, 3, 4, 6, 5, 5, 2, 3, 3, 1, 2, 5, 3, 7, 8, 4, 2, 3, 3, 2, 4, 1, 5, 1, 2, 2, 1, 3, 2, 2, 3, 3, 1, 4, 6, 1, 7, 2, 2, 3, 2, 4, 2, 2, 6, 1, 9, 3, 3, 3, 2, 2, 7, 3, 2, 5, 5, 4, 2, 2, 1, 6, 5, 9, 5, 3, 4, 5, 2, 4, 4, 3, 3, 2, 4, 4, 2, 1, 3, 4, 2, 2, 2, 4, 3, 2, 2, 5, 3, 8, 5, 4, 5, 1, 5, 3, 4, 1, 2, 3, 3, 8, 3, 2, 4, 4, 3, 3, 4, 6, 2, 4, 3, 2, 2, 8, 5, 2, 4, 2, 2, 2, 2, 4, 2, 6, 2, 2, 1, 2, 2, 4, 2, 3, 1, 7, 8, 2, 3, 5, 2, 2, 2, 2, 5, 4, 2, 4, 3, 3, 2, 3, 2, 2, 2, 2, 2, 3, 3, 3, 2 };
        @(posedge clk);
        val = '{ 2, 5, 4, 3, 3, 4, 3, 3, 7, 4, 5, 3, 5, 2, 1, 3, 3, 2, 9, 2, 2, 3, 4, 2, 1, 1, 3, 7, 4, 2, 3, 4, 2, 3, 3, 3, 2, 2, 3, 4, 2, 6, 3, 3, 5, 3, 3, 2, 2, 1, 3, 2, 8, 1, 2, 2, 4, 4, 2, 5, 2, 3, 4, 3, 3, 2, 4, 2, 2, 2, 6, 4, 2, 6, 6, 7, 3, 2, 4, 2, 4, 2, 2, 8, 6, 8, 6, 6, 2, 2, 5, 3, 3, 3, 7, 6, 2, 4, 3, 3, 3, 5, 5, 5, 3, 6, 5, 2, 3, 5, 1, 3, 1, 2, 5, 2, 2, 3, 5, 2, 2, 1, 6, 1, 4, 2, 6, 8, 3, 4, 3, 2, 4, 3, 4, 3, 2, 3, 3, 6, 1, 4, 2, 3, 4, 2, 2, 3, 5, 2, 4, 6, 1, 2, 1, 3, 3, 1, 1, 2, 2, 1, 3, 2, 8, 3, 2, 4, 2, 5, 6, 2, 7, 5, 9, 9, 2, 5, 2, 2, 4, 3, 3, 4, 3, 2, 4, 7, 2, 2, 2, 3, 2, 1, 2, 5, 6, 3, 2, 4 };
        @(posedge clk);
        val = '{ 2, 4, 4, 2, 4, 3, 4, 5, 6, 4, 4, 5, 2, 2, 4, 2, 3, 2, 6, 2, 1, 3, 4, 2, 4, 5, 9, 7, 7, 2, 2, 2, 3, 3, 1, 3, 2, 2, 3, 5, 2, 5, 4, 8, 5, 2, 3, 1, 3, 1, 3, 1, 2, 4, 2, 2, 1, 2, 7, 3, 6, 2, 2, 8, 3, 1, 3, 2, 2, 2, 6, 3, 2, 5, 4, 3, 5, 1, 4, 4, 6, 2, 4, 5, 3, 2, 5, 4, 3, 3, 3, 3, 4, 4, 2, 1, 2, 1, 3, 3, 9, 5, 6, 2, 3, 4, 6, 2, 1, 5, 3, 1, 2, 3, 2, 2, 3, 6, 5, 4, 2, 3, 1, 2, 5, 3, 3, 4, 7, 3, 4, 3, 4, 3, 4, 3, 3, 4, 2, 7, 2, 3, 1, 4, 1, 2, 3, 2, 2, 2, 3, 5, 2, 2, 2, 5, 1, 2, 1, 6, 3, 1, 4, 2, 5, 2, 2, 5, 2, 3, 5, 3, 4, 6, 9, 7, 2, 4, 3, 2, 2, 2, 2, 9, 6, 2, 3, 3, 2, 3, 6, 5, 2, 1, 2, 8, 4, 4, 3, 4 };
        @(posedge clk);
        val = '{ 3, 4, 4, 3, 4, 5, 4, 5, 4, 4, 5, 3, 2, 2, 3, 3, 1, 3, 5, 2, 2, 3, 7, 2, 2, 2, 3, 8, 4, 2, 2, 3, 1, 2, 2, 1, 4, 2, 2, 8, 2, 7, 4, 3, 6, 5, 3, 2, 3, 2, 4, 2, 6, 4, 3, 2, 3, 2, 1, 4, 1, 3, 5, 9, 2, 2, 5, 4, 2, 3, 2, 1, 5, 5, 7, 1, 2, 2, 4, 4, 3, 2, 2, 6, 4, 3, 3, 6, 2, 2, 4, 3, 3, 2, 3, 6, 2, 4, 9, 3, 6, 5, 4, 5, 3, 4, 3, 6, 5, 3, 4, 3, 2, 2, 2, 2, 5, 5, 4, 2, 5, 1, 4, 2, 2, 5, 5, 6, 3, 2, 3, 3, 2, 3, 2, 3, 2, 3, 3, 3, 3, 2, 4, 2, 2, 2, 2, 3, 3, 2, 5, 6, 6, 1, 3, 3, 1, 3, 2, 4, 1, 2, 3, 2, 6, 2, 6, 5, 6, 4, 1, 4, 4, 1, 6, 4, 2, 3, 2, 1, 1, 2, 2, 4, 6, 2, 1, 8, 4, 2, 1, 5, 2, 2, 2, 4, 2, 3, 3, 4 };
        @(posedge clk);
        val = '{ 4, 4, 4, 2, 2, 5, 2, 5, 6, 3, 4, 6, 2, 4, 2, 3, 2, 6, 3, 2, 4, 2, 4, 3, 1, 7, 2, 5, 6, 2, 2, 3, 4, 4, 1, 6, 2, 2, 3, 3, 2, 6, 2, 4, 2, 3, 3, 4, 1, 2, 5, 2, 6, 5, 3, 1, 3, 3, 4, 5, 3, 2, 2, 7, 2, 2, 4, 5, 2, 4, 2, 4, 2, 4, 4, 3, 3, 2, 4, 3, 4, 2, 2, 5, 3, 3, 7, 4, 1, 2, 2, 3, 5, 2, 2, 5, 2, 5, 2, 2, 5, 5, 2, 2, 3, 5, 6, 2, 3, 3, 2, 3, 2, 2, 3, 1, 5, 2, 2, 4, 4, 2, 4, 1, 2, 4, 6, 6, 5, 4, 5, 4, 5, 6, 2, 3, 2, 3, 4, 4, 3, 3, 4, 3, 2, 3, 3, 2, 3, 4, 3, 7, 4, 3, 4, 3, 4, 2, 1, 2, 3, 2, 2, 2, 2, 2, 3, 8, 1, 3, 8, 2, 3, 6, 3, 3, 2, 4, 3, 8, 2, 2, 1, 3, 5, 2, 1, 5, 2, 3, 6, 3, 2, 2, 2, 5, 3, 2, 2, 3 };
        @(posedge clk);
        val = '{ 5, 4, 3, 1, 3, 3, 3, 2, 4, 3, 4, 6, 2, 2, 2, 3, 3, 4, 4, 2, 3, 2, 3, 2, 3, 2, 3, 7, 3, 2, 2, 4, 3, 3, 2, 3, 2, 5, 2, 3, 2, 6, 5, 2, 3, 4, 8, 3, 2, 2, 4, 2, 5, 2, 2, 2, 2, 2, 5, 5, 4, 3, 2, 4, 2, 2, 4, 5, 4, 2, 6, 4, 3, 8, 2, 5, 4, 2, 2, 3, 5, 3, 3, 6, 2, 9, 3, 4, 2, 2, 2, 3, 3, 4, 4, 3, 3, 8, 2, 5, 2, 8, 5, 3, 3, 4, 5, 5, 4, 4, 3, 3, 2, 2, 3, 5, 5, 4, 6, 3, 3, 3, 2, 2, 3, 2, 9, 2, 3, 4, 7, 2, 2, 8, 3, 4, 2, 4, 2, 6, 3, 2, 1, 6, 5, 2, 2, 2, 5, 2, 2, 4, 1, 4, 5, 3, 2, 3, 1, 2, 3, 2, 2, 3, 2, 2, 4, 3, 2, 6, 2, 2, 3, 5, 5, 9, 6, 4, 4, 2, 2, 3, 4, 2, 3, 2, 3, 3, 3, 5, 4, 4, 1, 2, 1, 4, 6, 3, 2, 3 };
        @(posedge clk);
        val = '{ 3, 4, 3, 2, 3, 6, 6, 2, 9, 3, 4, 3, 2, 2, 2, 3, 2, 2, 7, 3, 2, 2, 2, 3, 3, 4, 3, 7, 4, 2, 1, 4, 4, 4, 2, 6, 4, 6, 5, 3, 3, 4, 3, 2, 3, 3, 3, 2, 2, 2, 6, 2, 2, 2, 2, 2, 3, 2, 2, 5, 3, 3, 5, 6, 3, 2, 6, 2, 4, 3, 5, 4, 2, 5, 4, 6, 1, 2, 4, 3, 4, 1, 3, 5, 6, 2, 3, 4, 3, 3, 2, 3, 4, 5, 4, 7, 1, 4, 3, 2, 2, 4, 3, 3, 3, 3, 7, 2, 3, 4, 2, 3, 4, 1, 3, 2, 3, 5, 4, 4, 4, 3, 1, 2, 5, 4, 6, 5, 9, 3, 7, 2, 5, 2, 3, 3, 2, 2, 5, 6, 8, 4, 2, 4, 4, 2, 1, 4, 3, 8, 3, 4, 4, 5, 2, 6, 2, 2, 2, 1, 2, 1, 4, 2, 2, 3, 3, 3, 2, 5, 4, 3, 3, 3, 4, 3, 2, 4, 4, 3, 2, 2, 1, 6, 5, 1, 2, 6, 3, 2, 5, 4, 2, 2, 1, 7, 5, 2, 3, 3 };
        @(posedge clk);
        val = '{ 4, 4, 2, 2, 5, 2, 4, 2, 6, 2, 4, 5, 2, 2, 5, 3, 3, 3, 3, 2, 3, 3, 4, 3, 3, 5, 4, 9, 5, 2, 2, 3, 2, 2, 2, 2, 5, 3, 2, 5, 2, 5, 4, 2, 1, 2, 5, 4, 2, 2, 3, 4, 4, 3, 3, 3, 3, 1, 2, 5, 4, 4, 5, 5, 2, 2, 9, 3, 1, 3, 4, 4, 6, 7, 5, 7, 2, 2, 5, 3, 4, 2, 2, 5, 5, 3, 7, 6, 3, 3, 2, 6, 2, 2, 4, 1, 6, 4, 3, 2, 2, 5, 2, 3, 1, 3, 5, 2, 2, 7, 5, 6, 8, 2, 3, 3, 5, 6, 4, 2, 4, 2, 2, 2, 2, 2, 4, 7, 8, 2, 3, 5, 1, 5, 3, 3, 3, 3, 2, 4, 2, 3, 2, 4, 2, 2, 2, 2, 5, 2, 4, 1, 2, 4, 7, 5, 2, 1, 8, 2, 4, 2, 2, 2, 9, 3, 3, 5, 1, 4, 3, 1, 5, 2, 7, 5, 2, 1, 2, 2, 2, 1, 2, 7, 5, 1, 2, 4, 5, 3, 3, 4, 2, 2, 2, 5, 3, 5, 3, 2 };
        @(posedge clk);
        val = '{ 5, 3, 4, 4, 3, 3, 3, 4, 9, 3, 4, 4, 2, 4, 7, 1, 3, 2, 5, 2, 2, 3, 5, 4, 3, 5, 8, 4, 4, 1, 2, 6, 5, 3, 1, 4, 2, 1, 5, 7, 3, 7, 4, 2, 5, 4, 5, 4, 2, 1, 3, 2, 4, 3, 3, 2, 3, 2, 3, 3, 2, 2, 3, 6, 3, 6, 4, 3, 2, 3, 6, 3, 2, 2, 7, 7, 3, 2, 2, 2, 2, 2, 2, 5, 2, 2, 6, 7, 3, 5, 6, 7, 3, 3, 3, 2, 2, 5, 5, 3, 2, 8, 3, 4, 5, 3, 6, 4, 5, 5, 3, 2, 5, 2, 3, 2, 2, 3, 2, 2, 2, 2, 7, 2, 4, 5, 4, 9, 8, 4, 5, 4, 3, 3, 2, 2, 2, 5, 3, 2, 3, 3, 4, 5, 2, 2, 1, 2, 5, 2, 5, 6, 3, 2, 1, 7, 3, 4, 3, 2, 1, 2, 4, 3, 7, 2, 4, 7, 2, 7, 5, 2, 8, 6, 4, 9, 1, 4, 4, 2, 2, 2, 6, 4, 3, 2, 1, 3, 3, 5, 2, 2, 5, 2, 2, 2, 5, 3, 7, 2 };
        @(posedge clk);
        val = '{ 3, 5, 3, 2, 1, 7, 3, 3, 4, 4, 4, 5, 2, 4, 2, 3, 2, 2, 4, 2, 2, 2, 2, 3, 1, 3, 2, 1, 4, 2, 4, 1, 2, 2, 3, 5, 3, 2, 5, 7, 2, 5, 4, 3, 4, 2, 5, 2, 6, 2, 7, 2, 7, 8, 2, 2, 5, 2, 6, 4, 3, 4, 3, 9, 3, 2, 9, 4, 2, 3, 3, 2, 3, 7, 7, 5, 4, 1, 2, 3, 4, 2, 2, 8, 4, 4, 4, 3, 3, 2, 8, 8, 4, 2, 8, 2, 3, 5, 5, 2, 5, 5, 7, 2, 4, 3, 7, 3, 5, 3, 3, 3, 2, 2, 3, 6, 5, 1, 6, 3, 4, 2, 4, 6, 2, 3, 4, 6, 8, 5, 3, 2, 2, 4, 4, 3, 2, 3, 3, 4, 5, 3, 2, 3, 9, 2, 2, 4, 9, 2, 4, 3, 4, 4, 3, 4, 4, 3, 5, 2, 2, 3, 4, 2, 7, 3, 3, 3, 2, 5, 4, 3, 2, 4, 8, 8, 1, 3, 1, 2, 2, 2, 6, 1, 8, 2, 1, 3, 1, 3, 6, 3, 2, 3, 2, 6, 6, 3, 2, 2 };
        @(posedge clk);
        val = '{ 2, 7, 3, 3, 1, 5, 4, 1, 4, 2, 5, 3, 1, 5, 7, 3, 3, 4, 4, 2, 2, 2, 3, 2, 2, 8, 4, 6, 4, 2, 1, 7, 4, 5, 2, 6, 2, 2, 8, 9, 4, 6, 7, 7, 4, 2, 3, 2, 2, 2, 6, 2, 7, 4, 2, 1, 2, 2, 5, 2, 4, 4, 4, 5, 1, 2, 2, 2, 6, 3, 4, 3, 5, 5, 2, 7, 3, 6, 3, 6, 3, 2, 2, 5, 4, 2, 3, 3, 2, 1, 7, 3, 2, 4, 4, 4, 2, 5, 8, 4, 2, 6, 4, 2, 5, 3, 6, 3, 2, 7, 6, 3, 3, 4, 3, 2, 2, 3, 3, 5, 5, 3, 6, 2, 4, 2, 4, 6, 4, 5, 2, 4, 2, 6, 3, 3, 2, 2, 2, 5, 4, 3, 2, 4, 3, 5, 3, 3, 8, 4, 3, 3, 2, 2, 7, 6, 2, 5, 5, 1, 3, 2, 4, 1, 6, 2, 3, 4, 2, 3, 2, 2, 9, 7, 5, 5, 4, 4, 2, 1, 7, 3, 2, 3, 2, 1, 2, 6, 3, 2, 5, 4, 1, 2, 2, 7, 5, 5, 1, 1 };
        @(posedge clk);
        val = '{ 2, 6, 3, 2, 5, 7, 3, 2, 5, 4, 5, 1, 2, 1, 2, 3, 4, 2, 6, 2, 2, 3, 5, 1, 3, 1, 8, 4, 4, 1, 1, 2, 2, 4, 4, 3, 2, 2, 8, 4, 3, 6, 5, 3, 4, 2, 3, 2, 5, 2, 2, 2, 7, 2, 4, 2, 2, 2, 2, 2, 3, 5, 5, 4, 2, 2, 6, 2, 1, 3, 3, 3, 1, 2, 2, 3, 5, 2, 4, 2, 4, 3, 4, 6, 6, 3, 4, 3, 2, 2, 3, 3, 4, 2, 4, 7, 3, 5, 2, 3, 3, 4, 3, 4, 1, 4, 4, 5, 3, 3, 3, 3, 4, 1, 3, 4, 5, 2, 4, 2, 5, 2, 1, 2, 4, 3, 5, 2, 8, 2, 5, 5, 1, 2, 5, 3, 2, 4, 2, 6, 2, 3, 1, 4, 3, 2, 3, 3, 3, 2, 3, 6, 6, 4, 6, 7, 2, 5, 4, 5, 2, 2, 4, 3, 7, 3, 3, 6, 2, 4, 2, 6, 3, 8, 4, 4, 3, 3, 2, 3, 2, 3, 2, 7, 7, 1, 2, 2, 1, 3, 6, 3, 1, 2, 2, 6, 2, 7, 2, 2 };
        @(posedge clk);
        val = '{ 2, 4, 4, 2, 2, 5, 4, 3, 6, 4, 3, 2, 2, 4, 6, 1, 2, 6, 5, 2, 3, 9, 3, 2, 2, 2, 9, 5, 5, 2, 2, 4, 3, 5, 3, 3, 5, 4, 5, 3, 3, 6, 5, 9, 9, 4, 4, 5, 2, 2, 3, 2, 8, 6, 2, 2, 1, 2, 3, 5, 3, 8, 3, 3, 3, 2, 7, 5, 6, 5, 3, 3, 1, 5, 9, 6, 2, 2, 2, 3, 3, 1, 2, 5, 6, 4, 7, 4, 2, 3, 2, 5, 4, 3, 3, 7, 4, 3, 2, 2, 2, 7, 3, 1, 3, 3, 5, 2, 2, 8, 2, 3, 1, 4, 3, 1, 3, 4, 2, 4, 3, 2, 4, 1, 5, 2, 3, 2, 8, 2, 2, 1, 3, 3, 3, 2, 2, 4, 3, 6, 3, 3, 1, 2, 2, 3, 2, 1, 3, 2, 4, 4, 8, 7, 7, 6, 3, 4, 3, 1, 2, 2, 3, 3, 2, 3, 5, 5, 2, 2, 3, 2, 4, 3, 7, 8, 1, 3, 4, 2, 6, 2, 5, 2, 3, 2, 5, 4, 3, 2, 5, 4, 2, 1, 2, 6, 2, 3, 2, 5 };
        @(posedge clk);
        val = '{ 2, 4, 1, 2, 2, 4, 5, 4, 3, 3, 5, 5, 2, 3, 9, 3, 3, 3, 4, 2, 2, 1, 3, 2, 2, 3, 4, 8, 4, 4, 1, 4, 4, 2, 2, 3, 2, 2, 2, 7, 2, 6, 6, 3, 4, 3, 2, 6, 5, 2, 5, 3, 4, 6, 2, 2, 3, 2, 6, 1, 3, 3, 3, 4, 2, 2, 7, 5, 2, 3, 7, 1, 1, 7, 5, 5, 2, 2, 3, 3, 5, 2, 3, 7, 6, 3, 2, 3, 6, 3, 7, 6, 4, 2, 1, 1, 4, 8, 4, 1, 5, 5, 6, 6, 2, 2, 5, 4, 3, 9, 2, 3, 2, 1, 2, 2, 3, 4, 6, 5, 3, 3, 3, 2, 5, 2, 3, 5, 6, 3, 4, 1, 4, 2, 4, 3, 2, 2, 3, 4, 7, 3, 9, 4, 4, 2, 1, 2, 5, 2, 4, 3, 7, 6, 5, 9, 2, 5, 2, 4, 3, 2, 3, 1, 7, 3, 3, 5, 1, 4, 2, 2, 4, 3, 6, 5, 2, 4, 3, 3, 3, 2, 5, 6, 5, 2, 2, 4, 3, 3, 6, 4, 2, 3, 2, 1, 3, 4, 5, 4 };
        @(posedge clk);
        val = '{ 2, 4, 2, 2, 2, 4, 6, 2, 1, 4, 4, 5, 2, 9, 2, 3, 3, 1, 5, 2, 2, 2, 9, 2, 5, 2, 2, 7, 4, 2, 2, 4, 2, 5, 2, 4, 3, 2, 3, 4, 2, 5, 5, 1, 3, 3, 2, 5, 2, 2, 3, 2, 6, 7, 2, 2, 2, 2, 2, 1, 4, 9, 1, 4, 2, 2, 4, 5, 3, 5, 6, 4, 2, 4, 4, 6, 6, 3, 3, 2, 2, 2, 2, 6, 3, 3, 1, 3, 5, 2, 2, 2, 4, 3, 5, 2, 2, 8, 6, 2, 3, 3, 3, 6, 2, 1, 9, 2, 2, 2, 2, 3, 2, 2, 2, 4, 5, 4, 6, 5, 3, 3, 3, 4, 5, 3, 3, 5, 9, 5, 6, 7, 1, 2, 3, 3, 1, 4, 1, 3, 6, 3, 3, 3, 3, 2, 2, 2, 7, 3, 3, 3, 3, 4, 7, 6, 2, 3, 1, 2, 2, 2, 2, 2, 4, 3, 5, 6, 2, 4, 2, 2, 6, 4, 5, 5, 2, 7, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 4, 3, 3, 2, 2, 1, 1, 2, 3, 8, 4 };
        @(posedge clk);
        val = '{ 2, 4, 2, 3, 3, 5, 3, 1, 9, 4, 3, 2, 2, 1, 6, 2, 2, 2, 6, 1, 2, 3, 2, 3, 2, 2, 7, 4, 3, 2, 2, 4, 2, 2, 5, 3, 1, 4, 2, 6, 3, 5, 3, 7, 4, 4, 3, 2, 3, 4, 6, 1, 9, 2, 3, 2, 5, 2, 6, 4, 2, 7, 2, 7, 2, 1, 7, 9, 3, 4, 2, 2, 2, 5, 2, 5, 3, 1, 3, 5, 3, 3, 4, 5, 2, 2, 6, 5, 8, 1, 5, 8, 4, 2, 1, 5, 6, 4, 3, 1, 4, 4, 4, 3, 3, 4, 5, 1, 2, 2, 6, 2, 2, 1, 3, 2, 3, 4, 3, 3, 4, 4, 7, 1, 2, 3, 6, 5, 7, 3, 4, 6, 5, 3, 2, 2, 1, 5, 3, 9, 4, 3, 1, 2, 2, 1, 1, 3, 2, 2, 6, 6, 3, 2, 2, 1, 2, 5, 4, 9, 2, 2, 4, 2, 7, 3, 3, 1, 2, 5, 8, 2, 6, 4, 6, 6, 3, 3, 3, 1, 3, 1, 1, 3, 9, 4, 3, 4, 3, 2, 6, 4, 2, 2, 3, 8, 3, 3, 2, 3 };
        @(posedge clk);
        val = '{ 2, 5, 3, 2, 3, 5, 5, 4, 7, 1, 4, 5, 2, 3, 7, 1, 3, 2, 6, 2, 2, 3, 3, 2, 3, 3, 4, 5, 8, 2, 2, 3, 4, 3, 7, 4, 2, 2, 2, 4, 4, 6, 6, 3, 2, 3, 3, 2, 2, 2, 6, 2, 3, 6, 6, 2, 1, 3, 2, 3, 2, 2, 2, 3, 2, 2, 5, 6, 5, 3, 7, 4, 2, 5, 4, 8, 1, 2, 2, 1, 2, 2, 2, 7, 5, 3, 6, 6, 3, 2, 2, 9, 4, 2, 3, 7, 2, 5, 1, 2, 6, 8, 2, 5, 2, 5, 9, 3, 3, 8, 2, 2, 1, 4, 3, 3, 4, 4, 2, 7, 4, 4, 2, 2, 7, 2, 6, 6, 1, 3, 3, 2, 2, 2, 4, 2, 3, 2, 2, 1, 3, 2, 8, 4, 6, 4, 2, 2, 4, 2, 3, 6, 7, 2, 5, 3, 3, 1, 4, 3, 2, 2, 5, 1, 7, 3, 3, 4, 1, 3, 2, 5, 4, 6, 4, 7, 3, 4, 4, 2, 2, 2, 2, 3, 3, 2, 1, 9, 2, 3, 3, 5, 4, 2, 2, 2, 2, 3, 7, 4 };
        @(posedge clk);
        val = '{ 8, 8, 4, 2, 2, 2, 3, 6, 4, 3, 4, 4, 2, 3, 8, 3, 3, 2, 4, 1, 2, 1, 4, 3, 2, 2, 7, 2, 5, 5, 2, 2, 4, 5, 2, 3, 1, 3, 3, 9, 2, 3, 7, 6, 5, 4, 5, 3, 5, 1, 8, 1, 9, 4, 3, 2, 2, 5, 6, 5, 4, 4, 4, 3, 3, 6, 1, 4, 5, 3, 2, 4, 5, 4, 3, 7, 3, 2, 2, 5, 2, 3, 3, 4, 5, 2, 3, 3, 3, 2, 2, 3, 4, 1, 5, 3, 4, 3, 4, 3, 3, 5, 7, 6, 3, 4, 3, 5, 2, 7, 3, 4, 3, 2, 4, 3, 3, 2, 4, 2, 4, 3, 7, 1, 6, 4, 5, 4, 7, 3, 5, 5, 3, 3, 2, 2, 2, 4, 8, 3, 6, 3, 8, 5, 3, 2, 2, 4, 9, 2, 3, 5, 4, 2, 5, 6, 6, 5, 6, 3, 3, 2, 3, 2, 4, 2, 1, 5, 2, 5, 8, 2, 5, 7, 7, 8, 2, 4, 2, 2, 1, 2, 2, 3, 5, 4, 3, 4, 3, 3, 4, 4, 2, 2, 2, 2, 2, 4, 2, 2 };
        @(posedge clk);
        val = '{ 2, 4, 3, 3, 3, 5, 3, 2, 7, 4, 5, 4, 2, 4, 7, 3, 3, 2, 4, 3, 3, 6, 4, 3, 1, 2, 9, 7, 9, 2, 2, 2, 3, 2, 2, 3, 3, 4, 3, 8, 2, 4, 6, 3, 2, 2, 4, 5, 2, 2, 6, 4, 4, 4, 6, 2, 5, 6, 1, 5, 3, 8, 3, 3, 1, 2, 9, 5, 4, 7, 4, 2, 3, 5, 7, 8, 4, 2, 4, 4, 5, 1, 2, 8, 5, 8, 6, 5, 5, 4, 1, 3, 3, 5, 5, 4, 3, 5, 2, 3, 3, 8, 2, 2, 3, 4, 6, 2, 2, 8, 3, 3, 2, 2, 2, 3, 5, 4, 4, 3, 4, 3, 6, 4, 2, 2, 4, 3, 7, 3, 4, 6, 1, 4, 4, 3, 2, 3, 2, 6, 3, 2, 2, 6, 2, 2, 1, 2, 2, 1, 4, 3, 3, 1, 8, 3, 2, 5, 1, 7, 6, 2, 4, 8, 4, 2, 6, 4, 2, 3, 2, 2, 5, 6, 7, 5, 1, 3, 2, 2, 5, 4, 2, 5, 4, 2, 3, 3, 2, 3, 4, 4, 2, 2, 2, 3, 2, 1, 5, 4 };
        @(posedge clk);
        val = '{ 2, 4, 4, 3, 4, 4, 4, 5, 7, 2, 3, 4, 2, 2, 3, 3, 2, 2, 6, 6, 2, 3, 5, 2, 2, 4, 7, 5, 5, 3, 4, 4, 4, 2, 6, 3, 9, 1, 4, 6, 2, 5, 5, 2, 2, 2, 3, 3, 5, 2, 2, 2, 7, 5, 2, 2, 5, 2, 5, 4, 3, 7, 1, 6, 2, 1, 3, 7, 5, 7, 7, 4, 2, 3, 6, 6, 3, 2, 2, 2, 4, 3, 2, 8, 4, 5, 2, 5, 4, 3, 9, 4, 4, 6, 6, 4, 1, 5, 3, 4, 2, 5, 2, 4, 3, 3, 4, 4, 3, 6, 7, 3, 3, 4, 3, 6, 3, 4, 4, 7, 3, 2, 2, 1, 2, 2, 4, 5, 5, 4, 6, 6, 6, 3, 2, 4, 5, 4, 4, 2, 9, 3, 2, 4, 2, 3, 2, 7, 7, 2, 4, 5, 2, 2, 3, 3, 2, 4, 3, 2, 2, 2, 4, 1, 5, 3, 1, 3, 4, 6, 3, 2, 4, 5, 7, 7, 2, 3, 1, 2, 4, 7, 4, 3, 6, 2, 2, 4, 4, 3, 3, 4, 2, 2, 2, 2, 4, 5, 5, 4 };
        @(posedge clk);
        val = '{ 5, 2, 2, 4, 2, 2, 4, 2, 5, 3, 4, 3, 3, 6, 2, 4, 1, 2, 3, 1, 1, 4, 1, 1, 3, 1, 9, 2, 6, 1, 2, 3, 2, 2, 1, 3, 2, 1, 4, 2, 3, 9, 3, 4, 5, 6, 5, 3, 2, 2, 1, 2, 5, 2, 4, 2, 1, 2, 2, 5, 6, 3, 2, 5, 1, 3, 4, 3, 2, 3, 5, 3, 2, 6, 4, 3, 3, 2, 1, 5, 4, 4, 2, 9, 6, 2, 6, 3, 4, 2, 2, 1, 4, 5, 5, 3, 2, 7, 5, 1, 4, 5, 3, 4, 3, 4, 6, 1, 4, 5, 3, 1, 2, 4, 2, 2, 4, 2, 7, 3, 4, 1, 7, 2, 4, 2, 6, 7, 6, 3, 4, 2, 3, 5, 1, 3, 4, 4, 3, 4, 1, 3, 2, 2, 3, 2, 2, 2, 8, 1, 4, 2, 4, 2, 5, 3, 5, 6, 3, 1, 4, 4, 4, 3, 5, 3, 2, 5, 2, 3, 5, 1, 2, 6, 7, 6, 1, 6, 1, 2, 2, 2, 2, 7, 2, 1, 2, 4, 1, 4, 5, 1, 1, 2, 2, 6, 3, 3, 9, 4 };
        @(posedge clk);
        val = '{ 5, 4, 2, 2, 3, 4, 3, 5, 5, 4, 7, 3, 1, 5, 2, 3, 7, 4, 5, 2, 5, 3, 7, 3, 3, 6, 2, 1, 6, 1, 2, 5, 1, 9, 2, 4, 2, 2, 4, 4, 2, 3, 7, 2, 2, 4, 4, 4, 1, 2, 3, 2, 6, 5, 2, 2, 6, 2, 2, 2, 2, 1, 3, 5, 2, 2, 7, 4, 4, 7, 2, 4, 3, 6, 4, 4, 1, 2, 2, 3, 3, 2, 3, 3, 1, 2, 2, 4, 2, 2, 9, 3, 4, 5, 4, 2, 5, 3, 4, 2, 3, 3, 1, 4, 2, 5, 5, 4, 2, 7, 4, 3, 4, 2, 2, 3, 2, 8, 5, 1, 1, 1, 4, 1, 4, 2, 5, 6, 8, 4, 5, 2, 2, 6, 3, 3, 1, 5, 4, 2, 6, 7, 2, 5, 5, 4, 2, 2, 7, 5, 4, 5, 2, 2, 4, 2, 3, 3, 5, 4, 3, 4, 2, 3, 5, 4, 4, 5, 2, 4, 5, 1, 4, 6, 5, 5, 2, 3, 4, 3, 2, 2, 5, 7, 4, 1, 2, 3, 3, 3, 4, 2, 2, 2, 2, 6, 4, 3, 6, 3 };
        @(posedge clk);
        val = '{ 5, 5, 4, 4, 3, 7, 4, 2, 4, 4, 3, 5, 2, 1, 6, 3, 3, 2, 4, 2, 3, 2, 6, 3, 3, 4, 3, 5, 9, 2, 2, 4, 2, 4, 1, 2, 2, 2, 5, 3, 1, 6, 4, 3, 5, 2, 3, 2, 2, 2, 3, 3, 7, 1, 3, 2, 1, 2, 2, 4, 3, 1, 1, 6, 3, 2, 6, 5, 3, 3, 4, 4, 7, 8, 4, 7, 3, 2, 3, 3, 1, 3, 1, 4, 5, 3, 7, 2, 2, 3, 3, 7, 3, 1, 5, 8, 2, 3, 5, 2, 6, 5, 3, 2, 3, 3, 6, 3, 2, 4, 1, 3, 3, 2, 2, 5, 5, 4, 5, 4, 4, 2, 2, 4, 6, 4, 5, 7, 4, 4, 8, 2, 4, 7, 3, 2, 1, 1, 2, 5, 4, 4, 2, 2, 1, 3, 2, 2, 2, 4, 2, 3, 6, 2, 8, 5, 5, 3, 4, 2, 4, 2, 4, 1, 5, 3, 4, 4, 2, 2, 5, 5, 7, 6, 5, 9, 3, 4, 3, 3, 4, 5, 4, 3, 7, 2, 2, 4, 2, 6, 2, 3, 2, 2, 2, 5, 3, 3, 1, 3 };
        @(posedge clk);
        val = '{ 8, 5, 3, 4, 3, 3, 6, 9, 5, 4, 4, 5, 2, 2, 2, 1, 2, 4, 3, 2, 5, 3, 3, 2, 4, 2, 2, 4, 5, 2, 2, 4, 2, 2, 1, 3, 5, 7, 3, 8, 2, 4, 7, 6, 5, 6, 3, 2, 3, 2, 1, 2, 7, 2, 3, 2, 1, 2, 2, 3, 5, 3, 1, 8, 3, 2, 9, 8, 5, 4, 3, 4, 2, 6, 6, 4, 2, 2, 3, 3, 4, 1, 2, 4, 2, 2, 6, 2, 5, 3, 2, 4, 4, 2, 1, 8, 4, 5, 2, 3, 1, 3, 3, 5, 3, 4, 4, 3, 4, 8, 4, 3, 2, 4, 2, 5, 5, 4, 6, 3, 4, 2, 5, 2, 4, 2, 8, 3, 4, 3, 3, 6, 3, 3, 3, 4, 4, 6, 2, 8, 5, 3, 3, 3, 4, 5, 2, 2, 7, 2, 4, 6, 6, 4, 1, 4, 3, 2, 1, 3, 1, 2, 4, 2, 5, 4, 5, 8, 2, 3, 3, 3, 6, 5, 5, 2, 2, 3, 5, 2, 6, 2, 2, 5, 4, 2, 2, 3, 3, 3, 4, 2, 2, 2, 2, 8, 1, 2, 2, 3 };
        @(posedge clk);
        val = '{ 3, 3, 3, 4, 1, 2, 3, 3, 9, 2, 4, 2, 2, 2, 1, 2, 1, 2, 2, 1, 1, 3, 3, 1, 3, 2, 3, 4, 5, 2, 3, 5, 3, 2, 2, 4, 2, 2, 3, 8, 8, 7, 6, 7, 4, 5, 5, 3, 1, 2, 6, 2, 4, 2, 5, 2, 2, 1, 2, 2, 4, 3, 1, 6, 3, 2, 5, 5, 2, 3, 5, 4, 3, 4, 2, 8, 1, 1, 1, 6, 4, 2, 2, 9, 4, 4, 4, 6, 2, 2, 2, 2, 4, 4, 5, 8, 4, 5, 2, 3, 2, 5, 3, 2, 5, 3, 6, 2, 5, 9, 2, 2, 2, 4, 3, 3, 5, 4, 5, 4, 5, 3, 1, 2, 3, 3, 6, 5, 4, 4, 3, 5, 2, 4, 2, 2, 3, 2, 3, 7, 6, 3, 1, 1, 2, 2, 2, 2, 4, 2, 4, 5, 3, 2, 7, 2, 2, 5, 5, 8, 1, 2, 2, 5, 3, 4, 4, 2, 2, 2, 3, 3, 1, 6, 6, 6, 4, 4, 2, 4, 2, 2, 1, 6, 3, 1, 2, 3, 2, 3, 4, 1, 2, 3, 2, 6, 5, 3, 6, 1 };
        @(posedge clk);
        val = '{ 4, 2, 6, 2, 2, 3, 3, 2, 4, 4, 6, 4, 2, 1, 4, 3, 3, 4, 2, 1, 3, 3, 6, 2, 2, 4, 3, 2, 4, 2, 2, 4, 4, 1, 2, 3, 3, 4, 4, 9, 3, 3, 7, 4, 4, 3, 3, 2, 2, 2, 5, 2, 3, 7, 5, 2, 2, 2, 5, 5, 4, 6, 1, 6, 4, 2, 9, 9, 7, 3, 3, 4, 6, 5, 3, 5, 5, 1, 3, 3, 1, 1, 2, 5, 5, 5, 1, 3, 3, 1, 3, 6, 4, 5, 4, 4, 2, 5, 2, 3, 4, 5, 2, 2, 3, 4, 6, 4, 4, 4, 4, 4, 3, 1, 3, 4, 4, 4, 5, 2, 4, 3, 5, 5, 2, 5, 6, 3, 8, 6, 8, 6, 3, 3, 2, 2, 1, 3, 2, 1, 8, 4, 3, 4, 2, 5, 3, 2, 3, 3, 3, 4, 6, 2, 8, 3, 2, 4, 5, 9, 2, 1, 3, 2, 6, 4, 3, 6, 2, 2, 1, 2, 4, 6, 4, 7, 1, 1, 2, 4, 2, 1, 2, 3, 3, 2, 2, 6, 7, 3, 4, 2, 1, 1, 2, 5, 4, 1, 3, 3 };
        @(posedge clk);
        val = '{ 4, 6, 3, 2, 2, 6, 2, 6, 7, 4, 6, 2, 2, 5, 6, 3, 1, 2, 5, 2, 3, 1, 1, 2, 3, 3, 3, 8, 4, 2, 3, 4, 3, 3, 7, 5, 6, 4, 3, 8, 3, 6, 5, 4, 1, 2, 2, 2, 7, 2, 7, 3, 4, 3, 2, 1, 2, 2, 4, 3, 2, 4, 5, 6, 2, 2, 3, 1, 5, 3, 3, 4, 2, 5, 2, 3, 2, 1, 2, 3, 5, 2, 1, 5, 4, 1, 4, 3, 2, 2, 3, 9, 4, 3, 5, 4, 2, 4, 3, 2, 5, 4, 1, 5, 3, 4, 5, 2, 4, 4, 9, 3, 1, 7, 2, 8, 2, 3, 5, 3, 4, 3, 2, 7, 5, 1, 6, 6, 7, 6, 6, 4, 5, 3, 2, 3, 2, 1, 2, 5, 3, 2, 1, 2, 3, 3, 2, 3, 3, 3, 4, 4, 6, 5, 3, 8, 7, 3, 1, 5, 3, 2, 5, 2, 7, 3, 6, 5, 2, 3, 3, 3, 7, 7, 8, 5, 2, 4, 4, 2, 1, 3, 3, 5, 4, 2, 1, 4, 1, 3, 3, 3, 2, 2, 4, 7, 2, 3, 7, 2 };
        @(posedge clk);
        val = '{ 3, 3, 2, 3, 4, 6, 4, 6, 7, 4, 4, 6, 2, 3, 7, 3, 2, 3, 3, 2, 2, 3, 5, 1, 3, 2, 7, 5, 8, 2, 2, 4, 2, 2, 1, 2, 2, 2, 2, 6, 2, 4, 6, 2, 2, 2, 6, 4, 6, 3, 6, 1, 4, 2, 3, 3, 2, 5, 2, 3, 6, 4, 5, 5, 2, 2, 3, 4, 3, 1, 4, 1, 2, 2, 2, 7, 3, 3, 2, 3, 4, 4, 2, 4, 2, 2, 7, 3, 3, 2, 6, 7, 2, 3, 2, 5, 2, 9, 5, 2, 1, 7, 3, 5, 1, 4, 3, 4, 4, 3, 4, 3, 2, 1, 3, 2, 5, 3, 6, 4, 4, 3, 3, 1, 4, 3, 4, 3, 8, 5, 5, 5, 2, 4, 3, 3, 3, 3, 2, 4, 3, 3, 2, 2, 2, 2, 2, 3, 3, 2, 2, 3, 6, 3, 7, 7, 2, 5, 2, 8, 2, 2, 3, 2, 7, 3, 3, 5, 2, 6, 1, 4, 3, 6, 7, 9, 2, 2, 2, 2, 2, 2, 3, 2, 6, 2, 3, 5, 2, 3, 5, 2, 3, 2, 2, 4, 4, 2, 5, 4 };
        @(posedge clk);
        val = '{ 3, 5, 4, 3, 3, 4, 3, 6, 7, 3, 4, 3, 2, 2, 5, 3, 3, 4, 3, 2, 1, 8, 3, 3, 2, 2, 4, 4, 3, 4, 2, 2, 2, 1, 6, 5, 2, 3, 1, 5, 2, 5, 4, 7, 3, 2, 5, 3, 2, 2, 4, 3, 4, 4, 1, 2, 3, 3, 4, 5, 3, 3, 2, 6, 2, 2, 2, 6, 2, 2, 6, 2, 2, 7, 2, 7, 9, 2, 2, 2, 3, 2, 4, 5, 6, 5, 1, 4, 3, 4, 2, 2, 3, 5, 5, 2, 2, 8, 3, 1, 2, 5, 2, 2, 3, 4, 4, 2, 2, 8, 3, 5, 2, 2, 6, 3, 2, 7, 6, 5, 3, 2, 2, 2, 7, 2, 6, 4, 8, 4, 3, 4, 4, 3, 3, 1, 3, 6, 3, 2, 5, 4, 5, 6, 4, 3, 3, 3, 4, 2, 3, 2, 2, 5, 1, 5, 7, 3, 5, 3, 3, 3, 3, 4, 8, 4, 2, 6, 3, 3, 2, 4, 8, 3, 5, 8, 2, 3, 2, 2, 2, 5, 1, 3, 3, 2, 3, 7, 2, 3, 3, 2, 2, 2, 1, 4, 5, 4, 6, 1 };
        @(posedge clk);
        val = '{ 5, 3, 6, 2, 2, 4, 2, 2, 8, 2, 4, 5, 2, 6, 5, 4, 2, 2, 5, 2, 2, 2, 3, 3, 2, 2, 1, 2, 7, 2, 2, 3, 2, 3, 3, 6, 2, 2, 2, 6, 3, 5, 3, 3, 5, 6, 4, 4, 8, 2, 5, 1, 4, 4, 3, 2, 2, 2, 2, 2, 4, 3, 4, 3, 3, 2, 7, 5, 2, 3, 2, 1, 4, 5, 5, 5, 4, 2, 1, 3, 3, 1, 2, 9, 3, 2, 3, 4, 5, 3, 5, 3, 4, 4, 5, 8, 2, 4, 4, 3, 2, 4, 2, 6, 2, 6, 6, 2, 3, 9, 3, 3, 2, 2, 3, 5, 6, 2, 4, 2, 1, 3, 6, 2, 2, 2, 6, 5, 3, 5, 8, 2, 2, 1, 4, 2, 4, 4, 3, 6, 2, 3, 3, 4, 3, 2, 6, 2, 3, 2, 4, 3, 3, 2, 6, 5, 2, 5, 2, 3, 2, 5, 4, 2, 2, 1, 1, 4, 2, 2, 3, 2, 2, 8, 1, 3, 2, 4, 2, 2, 2, 2, 2, 5, 6, 4, 1, 7, 3, 3, 4, 3, 2, 2, 2, 4, 1, 2, 3, 3 };
        @(posedge clk);
        val = '{ 1, 4, 3, 1, 2, 5, 2, 2, 8, 5, 6, 6, 1, 2, 5, 4, 3, 1, 4, 1, 2, 4, 4, 2, 3, 6, 4, 3, 3, 1, 2, 3, 2, 5, 2, 3, 3, 3, 3, 7, 1, 6, 3, 7, 4, 3, 2, 5, 2, 1, 3, 2, 5, 4, 5, 2, 2, 2, 1, 3, 3, 5, 3, 7, 2, 2, 3, 5, 7, 2, 3, 1, 2, 3, 7, 3, 5, 2, 1, 3, 4, 2, 2, 9, 7, 4, 2, 3, 5, 2, 6, 2, 3, 2, 7, 7, 2, 2, 3, 1, 3, 4, 2, 3, 2, 3, 4, 3, 3, 5, 4, 3, 3, 2, 3, 2, 2, 3, 7, 3, 2, 2, 3, 2, 2, 2, 6, 6, 7, 3, 3, 3, 3, 1, 3, 3, 2, 3, 4, 7, 6, 1, 2, 2, 3, 2, 2, 3, 5, 4, 4, 2, 4, 2, 1, 3, 2, 2, 5, 4, 3, 2, 4, 2, 7, 3, 8, 4, 2, 5, 5, 3, 4, 6, 7, 9, 2, 4, 4, 2, 2, 5, 2, 2, 6, 2, 6, 4, 3, 2, 3, 4, 2, 4, 1, 6, 3, 1, 2, 5 };
        @(posedge clk);
        val = '{ 2, 6, 1, 3, 3, 3, 5, 1, 5, 2, 4, 4, 2, 4, 2, 2, 2, 2, 7, 1, 2, 3, 3, 2, 2, 2, 3, 3, 3, 2, 2, 4, 4, 2, 2, 3, 2, 2, 5, 8, 1, 7, 7, 2, 3, 2, 3, 2, 5, 2, 3, 2, 7, 2, 3, 3, 1, 2, 4, 3, 4, 3, 1, 7, 2, 2, 6, 5, 1, 3, 4, 2, 2, 3, 1, 4, 4, 2, 4, 3, 7, 3, 4, 5, 3, 3, 5, 2, 2, 3, 2, 9, 3, 2, 2, 3, 3, 2, 2, 2, 3, 4, 3, 3, 3, 6, 6, 2, 3, 1, 3, 2, 2, 4, 3, 2, 2, 3, 6, 2, 8, 1, 4, 2, 3, 2, 3, 6, 5, 2, 3, 3, 2, 6, 1, 3, 4, 5, 3, 6, 6, 3, 4, 5, 3, 2, 2, 1, 2, 1, 3, 6, 4, 3, 8, 7, 4, 1, 2, 7, 1, 1, 2, 2, 7, 4, 5, 5, 2, 6, 8, 2, 9, 3, 6, 9, 1, 3, 2, 2, 2, 2, 2, 5, 3, 3, 3, 3, 2, 3, 4, 1, 2, 2, 2, 6, 2, 2, 2, 3 };
        @(posedge clk);
        val = '{ 3, 5, 4, 3, 2, 3, 3, 1, 8, 4, 4, 5, 3, 4, 4, 6, 1, 2, 9, 3, 5, 2, 2, 2, 4, 2, 8, 2, 6, 2, 2, 2, 2, 2, 2, 4, 5, 2, 8, 8, 8, 5, 5, 2, 4, 2, 3, 2, 3, 2, 6, 2, 6, 2, 3, 2, 1, 2, 1, 1, 4, 5, 2, 8, 2, 2, 3, 9, 2, 6, 3, 3, 4, 3, 4, 3, 4, 2, 3, 3, 2, 2, 2, 9, 4, 3, 4, 3, 3, 4, 2, 3, 4, 5, 4, 6, 3, 5, 4, 3, 5, 6, 1, 2, 3, 3, 7, 4, 8, 4, 3, 3, 4, 2, 3, 6, 5, 4, 4, 4, 4, 3, 3, 1, 4, 4, 3, 6, 4, 4, 5, 3, 2, 3, 5, 4, 4, 4, 1, 7, 6, 3, 2, 6, 2, 3, 2, 2, 3, 2, 3, 5, 3, 4, 6, 4, 2, 2, 1, 7, 1, 2, 3, 2, 1, 1, 2, 5, 3, 6, 4, 3, 4, 4, 6, 7, 3, 4, 2, 2, 6, 1, 4, 2, 9, 2, 1, 4, 3, 3, 3, 3, 2, 1, 2, 6, 6, 3, 3, 3 };
        @(posedge clk);
        val = '{ 4, 1, 3, 2, 1, 5, 3, 7, 6, 1, 3, 5, 3, 2, 4, 3, 3, 2, 5, 2, 2, 3, 3, 2, 3, 3, 8, 7, 5, 2, 2, 3, 4, 2, 3, 4, 2, 2, 3, 5, 2, 5, 4, 2, 4, 5, 3, 2, 2, 3, 3, 2, 5, 2, 6, 2, 3, 2, 5, 5, 4, 2, 5, 8, 2, 3, 5, 2, 2, 3, 5, 3, 3, 7, 7, 4, 2, 2, 1, 3, 3, 2, 4, 6, 3, 2, 2, 5, 2, 3, 5, 7, 3, 2, 2, 6, 3, 5, 3, 2, 3, 7, 3, 2, 3, 4, 4, 5, 3, 2, 3, 3, 1, 4, 3, 5, 5, 5, 6, 5, 4, 2, 5, 2, 6, 3, 2, 5, 5, 4, 3, 1, 3, 8, 2, 3, 2, 2, 3, 7, 4, 3, 5, 4, 3, 5, 1, 2, 3, 2, 5, 2, 7, 5, 2, 4, 2, 3, 5, 2, 2, 2, 4, 2, 3, 3, 2, 3, 2, 3, 5, 3, 7, 6, 2, 8, 2, 7, 1, 2, 5, 2, 3, 3, 5, 1, 2, 6, 2, 4, 4, 3, 2, 1, 2, 2, 7, 2, 2, 6 };
        @(posedge clk);
        val = '{ 5, 3, 7, 2, 3, 1, 2, 3, 6, 4, 2, 2, 1, 2, 5, 4, 3, 2, 4, 1, 1, 3, 6, 2, 2, 5, 6, 5, 3, 3, 2, 4, 2, 3, 1, 3, 3, 2, 3, 6, 2, 5, 3, 6, 4, 1, 5, 2, 4, 2, 2, 3, 6, 3, 2, 3, 3, 2, 1, 4, 2, 5, 5, 6, 3, 2, 4, 5, 4, 8, 7, 1, 2, 5, 2, 5, 3, 9, 3, 3, 3, 2, 1, 9, 3, 2, 1, 4, 3, 3, 6, 7, 2, 2, 5, 5, 2, 5, 2, 2, 6, 7, 2, 4, 3, 4, 6, 4, 3, 8, 4, 2, 1, 2, 3, 4, 6, 5, 5, 2, 3, 2, 6, 2, 2, 3, 3, 4, 3, 3, 6, 3, 1, 1, 3, 3, 4, 4, 2, 5, 5, 3, 2, 4, 3, 2, 2, 2, 3, 2, 4, 1, 4, 4, 7, 5, 3, 4, 1, 2, 2, 2, 2, 2, 8, 6, 5, 5, 2, 7, 6, 2, 4, 5, 3, 6, 1, 2, 2, 2, 1, 3, 3, 2, 3, 2, 2, 5, 3, 7, 5, 2, 2, 2, 2, 7, 2, 3, 1, 2 };
        @(posedge clk);
        val = '{ 5, 4, 5, 2, 3, 5, 3, 3, 3, 3, 4, 1, 2, 2, 1, 3, 1, 2, 4, 2, 7, 3, 2, 2, 2, 1, 3, 5, 8, 2, 2, 1, 4, 2, 2, 4, 3, 1, 3, 6, 2, 6, 2, 9, 1, 6, 5, 2, 3, 2, 3, 1, 6, 3, 2, 2, 4, 5, 2, 2, 8, 2, 3, 3, 2, 2, 2, 4, 3, 5, 7, 3, 2, 5, 2, 4, 1, 5, 3, 2, 6, 2, 2, 5, 2, 3, 2, 1, 2, 3, 2, 8, 4, 3, 2, 2, 2, 5, 3, 3, 5, 5, 2, 5, 1, 3, 5, 5, 4, 7, 3, 4, 2, 4, 5, 2, 2, 4, 6, 3, 4, 1, 2, 3, 4, 2, 3, 6, 5, 6, 2, 3, 2, 3, 5, 4, 1, 5, 2, 1, 5, 3, 2, 2, 3, 2, 2, 2, 2, 2, 4, 6, 7, 3, 3, 4, 2, 5, 4, 8, 2, 2, 3, 2, 8, 4, 4, 5, 2, 3, 1, 6, 5, 9, 2, 9, 2, 3, 2, 1, 2, 2, 2, 2, 9, 2, 2, 3, 2, 4, 5, 2, 2, 2, 2, 3, 2, 5, 2, 2 };
        @(posedge clk);
        val = '{ 3, 6, 3, 2, 2, 4, 3, 3, 9, 4, 4, 5, 2, 2, 4, 3, 5, 2, 5, 2, 2, 6, 4, 3, 2, 2, 4, 5, 3, 1, 1, 4, 5, 2, 3, 4, 6, 2, 8, 5, 2, 6, 3, 6, 5, 3, 5, 4, 3, 2, 2, 2, 3, 3, 4, 2, 4, 2, 3, 3, 4, 2, 4, 2, 3, 2, 5, 3, 4, 3, 5, 1, 1, 3, 2, 5, 3, 2, 3, 7, 4, 2, 2, 5, 2, 2, 3, 3, 3, 2, 2, 5, 3, 2, 5, 2, 6, 2, 3, 3, 2, 4, 4, 5, 5, 4, 4, 2, 2, 7, 2, 3, 1, 4, 3, 6, 4, 8, 6, 1, 2, 1, 3, 2, 6, 2, 5, 6, 1, 3, 2, 4, 4, 5, 2, 3, 3, 5, 2, 3, 5, 2, 9, 6, 1, 2, 3, 1, 7, 3, 3, 1, 6, 6, 4, 6, 2, 2, 6, 1, 2, 2, 2, 3, 5, 3, 2, 7, 2, 3, 3, 2, 5, 5, 3, 9, 2, 3, 2, 2, 3, 2, 3, 3, 1, 1, 4, 1, 3, 4, 3, 5, 2, 2, 2, 6, 4, 3, 2, 4 };
        @(posedge clk);
        val = '{ 2, 6, 2, 2, 3, 4, 2, 7, 5, 4, 3, 5, 2, 2, 1, 3, 4, 2, 5, 2, 2, 3, 3, 2, 3, 4, 2, 6, 4, 3, 3, 2, 4, 3, 2, 3, 6, 5, 3, 5, 2, 4, 4, 6, 1, 2, 5, 3, 2, 1, 3, 4, 3, 3, 3, 2, 4, 2, 2, 3, 2, 4, 3, 1, 5, 2, 3, 2, 2, 3, 4, 3, 2, 4, 9, 9, 2, 2, 3, 4, 4, 5, 2, 6, 4, 2, 4, 4, 5, 3, 1, 4, 4, 5, 3, 6, 3, 5, 4, 2, 1, 5, 4, 3, 7, 5, 5, 4, 4, 7, 4, 3, 2, 4, 3, 3, 4, 2, 6, 5, 3, 3, 6, 1, 4, 1, 6, 4, 3, 5, 6, 1, 3, 6, 2, 4, 2, 4, 4, 3, 7, 1, 2, 2, 3, 2, 2, 2, 4, 4, 3, 1, 3, 3, 7, 4, 3, 3, 2, 5, 3, 3, 3, 2, 6, 3, 3, 5, 1, 3, 6, 2, 3, 2, 3, 9, 3, 3, 2, 2, 2, 5, 2, 1, 2, 2, 2, 5, 3, 5, 4, 4, 2, 1, 2, 6, 2, 3, 2, 4 };
        @(posedge clk);
        val = '{ 5, 5, 6, 1, 2, 3, 3, 5, 4, 5, 5, 5, 2, 1, 3, 4, 6, 2, 4, 1, 2, 5, 3, 2, 3, 3, 2, 7, 5, 4, 3, 4, 3, 4, 3, 8, 6, 2, 5, 3, 4, 3, 5, 4, 4, 2, 4, 8, 4, 2, 5, 2, 3, 2, 5, 2, 2, 2, 1, 2, 2, 3, 4, 5, 1, 2, 1, 2, 2, 4, 7, 4, 2, 7, 4, 8, 3, 4, 3, 3, 4, 2, 4, 8, 5, 4, 4, 7, 2, 3, 2, 2, 4, 2, 5, 2, 2, 5, 3, 1, 3, 5, 2, 5, 3, 4, 6, 7, 5, 8, 2, 3, 4, 3, 3, 2, 3, 3, 5, 1, 4, 2, 6, 2, 5, 2, 5, 5, 5, 4, 4, 7, 3, 5, 3, 3, 2, 7, 5, 4, 2, 2, 1, 2, 2, 4, 2, 1, 3, 2, 3, 5, 3, 3, 2, 3, 4, 3, 2, 3, 3, 1, 2, 2, 6, 3, 5, 5, 2, 3, 3, 3, 3, 2, 8, 6, 2, 4, 2, 1, 2, 2, 7, 7, 5, 2, 2, 2, 3, 3, 4, 2, 2, 2, 2, 5, 3, 3, 2, 1 };
        @(posedge clk);
        val = '{ 3, 5, 3, 3, 1, 5, 7, 1, 7, 3, 4, 2, 2, 6, 8, 5, 6, 1, 8, 2, 2, 5, 3, 2, 2, 4, 4, 4, 6, 2, 1, 1, 3, 4, 3, 1, 1, 2, 3, 8, 2, 5, 5, 5, 5, 2, 4, 3, 8, 3, 3, 2, 6, 2, 2, 2, 3, 4, 5, 2, 4, 3, 1, 6, 1, 2, 3, 9, 2, 5, 1, 4, 2, 6, 2, 7, 1, 2, 4, 4, 4, 5, 2, 6, 3, 3, 6, 4, 3, 3, 4, 8, 4, 3, 5, 7, 3, 2, 9, 7, 1, 3, 4, 4, 6, 3, 4, 5, 3, 8, 2, 3, 3, 4, 3, 1, 2, 4, 5, 4, 2, 3, 5, 2, 6, 4, 6, 7, 3, 7, 4, 2, 4, 5, 3, 3, 2, 3, 1, 3, 3, 7, 2, 6, 7, 3, 4, 3, 8, 2, 3, 6, 3, 2, 2, 4, 6, 5, 5, 3, 1, 2, 4, 2, 5, 3, 1, 4, 1, 6, 2, 2, 6, 9, 3, 7, 1, 3, 1, 1, 2, 2, 1, 4, 7, 2, 1, 7, 3, 3, 8, 2, 3, 4, 2, 2, 4, 5, 1, 5 };
        @(posedge clk);
        val = '{ 5, 4, 5, 2, 2, 2, 6, 3, 4, 2, 6, 5, 1, 5, 3, 3, 4, 2, 4, 6, 3, 2, 3, 2, 3, 2, 2, 9, 6, 4, 2, 5, 2, 3, 2, 6, 2, 1, 3, 4, 1, 4, 7, 3, 4, 3, 3, 4, 6, 2, 4, 2, 3, 7, 1, 2, 2, 2, 1, 2, 4, 3, 2, 4, 2, 2, 4, 7, 2, 2, 6, 1, 2, 6, 2, 2, 3, 3, 4, 3, 3, 2, 2, 5, 4, 3, 4, 6, 1, 1, 4, 3, 4, 2, 5, 2, 2, 5, 2, 3, 4, 6, 1, 5, 2, 5, 5, 1, 3, 2, 2, 5, 1, 2, 2, 1, 3, 4, 8, 1, 6, 2, 1, 2, 3, 4, 6, 5, 5, 7, 4, 3, 3, 2, 2, 3, 3, 3, 2, 2, 2, 6, 2, 3, 2, 3, 2, 1, 1, 4, 7, 3, 5, 2, 4, 5, 3, 6, 2, 2, 1, 2, 3, 2, 6, 1, 3, 5, 2, 2, 2, 3, 3, 5, 4, 6, 5, 8, 4, 2, 4, 5, 2, 3, 4, 4, 2, 4, 2, 5, 3, 1, 3, 2, 2, 5, 3, 3, 2, 3 };
        @(posedge clk);
        val = '{ 2, 7, 4, 2, 2, 5, 2, 2, 9, 4, 5, 5, 1, 2, 7, 2, 2, 2, 5, 2, 2, 3, 4, 2, 2, 4, 2, 5, 3, 4, 2, 2, 2, 2, 2, 4, 2, 2, 5, 5, 4, 6, 2, 3, 4, 3, 3, 2, 5, 2, 7, 2, 5, 6, 3, 2, 2, 2, 1, 2, 3, 3, 3, 1, 1, 2, 3, 3, 2, 3, 3, 1, 2, 5, 7, 8, 3, 2, 7, 5, 6, 2, 4, 9, 4, 4, 6, 5, 2, 3, 3, 6, 3, 2, 1, 3, 2, 4, 8, 3, 1, 6, 3, 2, 3, 2, 5, 2, 2, 6, 3, 4, 2, 1, 3, 1, 5, 2, 3, 5, 3, 4, 5, 2, 6, 2, 3, 5, 4, 2, 4, 2, 2, 2, 2, 5, 2, 4, 4, 6, 4, 3, 5, 2, 2, 2, 2, 2, 2, 2, 4, 5, 4, 4, 2, 7, 4, 3, 5, 2, 2, 2, 4, 1, 5, 2, 5, 7, 1, 3, 4, 2, 4, 3, 4, 6, 2, 2, 4, 4, 2, 2, 3, 6, 2, 4, 3, 4, 2, 2, 2, 4, 1, 1, 2, 5, 2, 3, 2, 4 };
        @(posedge clk);
        val = '{ 4, 4, 5, 2, 2, 7, 3, 4, 4, 3, 4, 1, 2, 4, 4, 2, 2, 4, 5, 2, 2, 2, 4, 2, 2, 5, 5, 8, 3, 3, 3, 1, 2, 1, 3, 4, 2, 2, 5, 7, 3, 4, 3, 3, 4, 5, 3, 2, 2, 2, 2, 2, 1, 3, 3, 2, 3, 2, 2, 5, 4, 3, 1, 4, 2, 3, 5, 5, 3, 4, 2, 4, 2, 5, 5, 6, 3, 3, 2, 5, 4, 1, 1, 8, 4, 4, 4, 4, 2, 2, 5, 6, 3, 2, 6, 5, 4, 5, 2, 3, 4, 3, 2, 3, 2, 5, 4, 5, 5, 9, 2, 3, 5, 3, 3, 5, 5, 4, 8, 3, 3, 2, 3, 2, 4, 5, 6, 4, 6, 4, 6, 4, 3, 5, 2, 3, 4, 4, 1, 6, 4, 2, 5, 4, 1, 2, 4, 2, 4, 1, 2, 4, 6, 4, 4, 7, 4, 6, 1, 3, 2, 2, 5, 3, 8, 3, 2, 4, 2, 3, 3, 4, 3, 5, 5, 4, 2, 3, 5, 2, 1, 3, 2, 5, 6, 1, 2, 2, 2, 2, 6, 3, 2, 3, 2, 3, 3, 2, 3, 1 };
        @(posedge clk);
        val = '{ 2, 4, 1, 3, 3, 5, 3, 2, 4, 4, 2, 4, 2, 2, 3, 3, 3, 3, 3, 3, 2, 3, 5, 3, 3, 5, 7, 7, 3, 2, 2, 2, 2, 4, 3, 5, 2, 2, 2, 5, 2, 7, 3, 3, 4, 1, 4, 1, 7, 2, 7, 2, 3, 5, 7, 3, 3, 3, 2, 2, 2, 4, 5, 4, 3, 5, 1, 4, 2, 3, 1, 3, 4, 4, 3, 8, 3, 2, 1, 3, 4, 2, 4, 9, 5, 2, 5, 3, 6, 1, 2, 6, 4, 4, 5, 2, 2, 5, 2, 2, 3, 5, 3, 5, 3, 2, 4, 5, 5, 2, 3, 3, 2, 4, 3, 2, 2, 8, 6, 5, 4, 2, 5, 2, 2, 4, 5, 5, 6, 5, 3, 5, 2, 3, 4, 3, 1, 4, 2, 4, 2, 3, 3, 3, 1, 2, 2, 2, 7, 2, 3, 3, 4, 2, 8, 2, 2, 1, 2, 8, 2, 2, 4, 3, 7, 4, 2, 2, 2, 5, 2, 2, 3, 5, 8, 5, 2, 4, 1, 3, 2, 2, 4, 3, 6, 3, 2, 3, 1, 2, 2, 3, 2, 2, 2, 3, 5, 4, 2, 4 };
        @(posedge clk);
        val = '{ 6, 7, 4, 1, 2, 3, 3, 2, 6, 3, 4, 6, 3, 5, 2, 3, 3, 2, 6, 2, 3, 3, 4, 1, 2, 1, 8, 6, 5, 2, 2, 2, 1, 2, 3, 4, 2, 2, 5, 3, 2, 4, 4, 3, 5, 2, 6, 2, 3, 2, 4, 3, 3, 3, 1, 2, 3, 2, 3, 9, 5, 3, 1, 7, 2, 1, 6, 7, 1, 3, 2, 2, 1, 5, 4, 3, 3, 2, 3, 4, 2, 4, 4, 8, 2, 3, 1, 3, 3, 2, 5, 2, 2, 2, 4, 6, 2, 5, 3, 3, 3, 5, 2, 4, 4, 4, 5, 1, 2, 4, 3, 7, 2, 2, 3, 2, 6, 2, 6, 4, 5, 1, 3, 6, 2, 2, 6, 9, 3, 4, 5, 4, 2, 1, 1, 2, 2, 4, 3, 4, 3, 3, 2, 3, 7, 7, 2, 3, 3, 4, 8, 4, 4, 2, 1, 2, 2, 1, 3, 4, 3, 2, 3, 5, 9, 2, 3, 6, 2, 4, 2, 5, 3, 6, 3, 8, 3, 7, 2, 2, 1, 1, 3, 3, 4, 1, 2, 9, 3, 5, 3, 4, 3, 2, 2, 6, 3, 7, 3, 3 };
        @(posedge clk);
        val = '{ 4, 3, 2, 3, 1, 5, 3, 2, 9, 4, 4, 4, 2, 3, 2, 2, 3, 2, 6, 5, 4, 2, 5, 1, 3, 5, 2, 5, 1, 2, 2, 3, 1, 5, 3, 4, 2, 2, 2, 5, 2, 2, 5, 2, 4, 2, 4, 4, 5, 2, 4, 2, 4, 8, 6, 1, 5, 2, 5, 5, 4, 3, 3, 5, 3, 2, 4, 4, 2, 3, 6, 2, 2, 8, 4, 3, 2, 2, 4, 3, 2, 3, 1, 9, 2, 6, 7, 4, 2, 2, 2, 6, 2, 3, 4, 7, 2, 5, 2, 1, 3, 5, 1, 4, 1, 4, 6, 1, 2, 5, 2, 2, 5, 2, 3, 2, 4, 4, 4, 3, 3, 2, 3, 1, 4, 2, 4, 4, 8, 5, 6, 5, 3, 6, 1, 4, 2, 4, 4, 6, 7, 4, 2, 2, 2, 2, 2, 5, 4, 4, 2, 2, 3, 5, 6, 4, 4, 3, 3, 3, 3, 2, 2, 1, 2, 3, 2, 6, 9, 3, 3, 1, 4, 6, 6, 5, 2, 3, 2, 1, 2, 3, 8, 6, 3, 2, 4, 4, 4, 3, 4, 3, 3, 3, 1, 3, 2, 3, 5, 2 };
        @(posedge clk);
        val = '{ 2, 4, 4, 2, 4, 3, 2, 2, 7, 4, 6, 5, 2, 2, 3, 4, 2, 3, 4, 2, 2, 1, 4, 2, 4, 2, 4, 8, 4, 2, 1, 5, 2, 3, 2, 2, 3, 2, 3, 9, 2, 6, 4, 5, 2, 2, 3, 3, 7, 2, 6, 2, 4, 6, 3, 2, 2, 2, 3, 1, 2, 3, 5, 4, 3, 2, 8, 5, 4, 4, 6, 2, 3, 5, 1, 8, 6, 2, 4, 5, 5, 2, 2, 9, 5, 4, 1, 3, 2, 1, 2, 2, 1, 2, 2, 8, 2, 4, 2, 3, 2, 6, 2, 4, 2, 3, 8, 1, 3, 4, 2, 3, 5, 2, 5, 7, 5, 3, 6, 2, 4, 1, 6, 2, 3, 4, 4, 6, 9, 5, 3, 4, 1, 4, 3, 3, 2, 5, 2, 4, 4, 6, 2, 5, 1, 2, 4, 1, 7, 3, 5, 1, 4, 3, 7, 6, 3, 2, 4, 8, 3, 1, 4, 2, 8, 3, 3, 4, 2, 1, 1, 3, 5, 3, 4, 3, 3, 2, 1, 2, 3, 2, 3, 3, 9, 2, 2, 6, 3, 3, 3, 5, 2, 5, 2, 2, 4, 3, 2, 4 };
        @(posedge clk);
        val = '{ 2, 2, 4, 3, 2, 3, 3, 5, 7, 4, 5, 6, 2, 6, 2, 5, 2, 2, 5, 1, 1, 2, 1, 3, 2, 2, 4, 2, 4, 1, 3, 4, 2, 4, 2, 3, 5, 7, 5, 5, 2, 7, 6, 8, 3, 2, 3, 3, 6, 2, 3, 4, 2, 5, 3, 2, 3, 2, 3, 8, 6, 6, 5, 5, 1, 4, 3, 6, 2, 1, 2, 2, 2, 3, 9, 3, 3, 1, 2, 2, 4, 2, 1, 8, 4, 2, 1, 3, 1, 4, 1, 7, 5, 2, 3, 4, 2, 5, 3, 2, 6, 5, 6, 2, 2, 2, 4, 5, 2, 5, 2, 4, 2, 4, 3, 4, 5, 1, 4, 3, 3, 2, 2, 2, 6, 3, 5, 6, 6, 4, 6, 3, 3, 3, 4, 3, 3, 7, 4, 2, 7, 7, 2, 3, 2, 2, 2, 1, 1, 2, 4, 5, 3, 2, 1, 4, 1, 1, 5, 5, 2, 2, 4, 2, 1, 4, 2, 7, 3, 3, 7, 4, 4, 6, 6, 6, 4, 4, 2, 2, 1, 2, 5, 2, 6, 3, 2, 4, 3, 3, 4, 3, 1, 2, 2, 6, 4, 3, 4, 3 };
        @(posedge clk);
        val = '{ 3, 5, 4, 3, 3, 3, 7, 4, 5, 3, 4, 1, 2, 2, 4, 4, 3, 2, 6, 2, 5, 3, 3, 3, 3, 2, 8, 5, 5, 1, 1, 1, 3, 2, 2, 6, 6, 1, 5, 4, 2, 5, 2, 3, 6, 2, 3, 4, 3, 2, 3, 2, 2, 6, 3, 2, 2, 2, 2, 3, 3, 1, 1, 5, 2, 2, 6, 4, 4, 3, 7, 1, 2, 7, 3, 6, 3, 2, 2, 2, 3, 2, 1, 6, 5, 3, 1, 2, 3, 3, 6, 9, 5, 1, 2, 3, 2, 4, 1, 3, 2, 6, 3, 5, 3, 4, 5, 2, 3, 5, 1, 3, 4, 2, 2, 4, 5, 1, 6, 2, 7, 3, 3, 2, 3, 4, 9, 3, 7, 6, 3, 3, 2, 1, 4, 3, 1, 3, 1, 5, 3, 4, 3, 3, 2, 4, 2, 1, 4, 3, 4, 4, 5, 4, 6, 1, 2, 4, 2, 2, 2, 2, 4, 2, 2, 3, 5, 8, 2, 2, 3, 4, 2, 3, 9, 7, 1, 1, 2, 2, 4, 2, 2, 5, 4, 2, 2, 4, 1, 4, 6, 3, 5, 2, 2, 4, 3, 2, 1, 2 };
        @(posedge clk);
        val = '{ 5, 7, 3, 3, 3, 3, 3, 6, 8, 4, 3, 1, 2, 2, 5, 3, 2, 3, 2, 3, 2, 1, 4, 2, 3, 1, 4, 7, 6, 3, 3, 4, 4, 2, 2, 1, 1, 2, 6, 4, 2, 6, 8, 7, 1, 2, 3, 3, 2, 1, 3, 2, 4, 4, 2, 1, 2, 5, 5, 4, 3, 4, 5, 5, 3, 2, 1, 9, 3, 4, 6, 1, 2, 2, 4, 3, 6, 2, 4, 3, 5, 2, 2, 7, 3, 2, 4, 4, 7, 1, 2, 3, 1, 5, 5, 7, 2, 5, 2, 1, 2, 6, 3, 1, 3, 4, 1, 2, 3, 9, 4, 3, 2, 1, 4, 2, 3, 4, 4, 2, 7, 2, 4, 2, 3, 3, 9, 5, 7, 7, 4, 2, 5, 7, 3, 4, 4, 6, 2, 2, 5, 2, 2, 3, 7, 3, 2, 2, 4, 1, 2, 5, 3, 7, 6, 3, 5, 5, 2, 6, 2, 1, 4, 2, 8, 1, 3, 4, 2, 1, 5, 4, 4, 3, 6, 6, 2, 3, 4, 8, 2, 2, 5, 2, 5, 3, 2, 3, 1, 2, 3, 4, 2, 2, 2, 7, 2, 2, 2, 3 };
        @(posedge clk);
        val = '{ 3, 4, 1, 5, 4, 5, 3, 2, 4, 5, 2, 3, 2, 2, 7, 4, 3, 6, 5, 2, 3, 5, 4, 2, 4, 2, 2, 5, 4, 2, 2, 2, 2, 2, 7, 4, 2, 7, 3, 4, 4, 5, 7, 3, 2, 2, 3, 1, 5, 2, 8, 1, 4, 3, 3, 2, 4, 2, 7, 8, 3, 8, 4, 9, 2, 2, 6, 5, 5, 4, 6, 1, 1, 3, 7, 6, 3, 2, 6, 5, 5, 2, 2, 9, 5, 2, 1, 5, 3, 3, 3, 1, 3, 2, 7, 3, 2, 9, 2, 3, 3, 5, 3, 2, 2, 1, 6, 1, 3, 6, 3, 1, 3, 1, 3, 7, 5, 6, 5, 2, 4, 2, 3, 2, 6, 3, 2, 4, 7, 4, 3, 1, 2, 7, 2, 3, 2, 6, 2, 1, 3, 3, 8, 3, 2, 3, 2, 2, 3, 2, 3, 2, 7, 4, 6, 3, 1, 6, 2, 4, 3, 3, 2, 4, 5, 3, 4, 4, 1, 4, 4, 2, 5, 7, 3, 6, 2, 3, 2, 2, 5, 5, 5, 3, 1, 1, 4, 3, 2, 3, 3, 3, 5, 1, 2, 6, 5, 3, 2, 2 };
        @(posedge clk);
        val = '{ 2, 6, 3, 3, 3, 4, 3, 4, 5, 3, 3, 5, 1, 4, 6, 2, 8, 3, 4, 2, 2, 5, 4, 2, 2, 5, 3, 6, 6, 2, 2, 2, 2, 2, 2, 4, 6, 4, 3, 4, 1, 9, 5, 3, 5, 2, 3, 4, 2, 2, 6, 2, 4, 5, 5, 1, 3, 2, 1, 3, 8, 3, 3, 7, 1, 2, 7, 5, 2, 5, 6, 4, 2, 1, 6, 9, 5, 5, 3, 4, 4, 3, 2, 8, 4, 3, 3, 4, 3, 3, 4, 7, 4, 1, 3, 4, 2, 4, 4, 2, 2, 5, 5, 4, 3, 3, 5, 5, 7, 8, 3, 3, 2, 2, 4, 2, 6, 7, 6, 4, 1, 3, 4, 2, 3, 2, 4, 8, 6, 6, 2, 4, 5, 2, 2, 2, 2, 5, 4, 3, 2, 3, 2, 4, 5, 3, 2, 2, 4, 2, 2, 5, 7, 3, 5, 2, 2, 1, 3, 6, 2, 2, 3, 2, 6, 3, 5, 5, 2, 3, 2, 2, 8, 2, 2, 6, 7, 3, 2, 2, 2, 1, 2, 3, 8, 1, 3, 4, 3, 3, 4, 3, 2, 2, 1, 4, 4, 2, 2, 4 };
        @(posedge clk);
        val = '{ 4, 4, 5, 2, 3, 5, 3, 2, 5, 3, 3, 4, 1, 1, 2, 4, 4, 3, 6, 2, 3, 3, 3, 3, 2, 4, 3, 3, 4, 2, 2, 3, 2, 2, 3, 4, 2, 2, 3, 5, 2, 3, 3, 3, 2, 4, 7, 2, 6, 2, 3, 2, 4, 2, 3, 3, 1, 4, 5, 2, 4, 7, 2, 3, 2, 2, 6, 4, 8, 4, 2, 3, 2, 7, 2, 3, 2, 2, 2, 2, 4, 2, 3, 7, 5, 3, 2, 4, 3, 2, 3, 8, 4, 1, 5, 2, 2, 4, 3, 2, 1, 5, 1, 3, 3, 5, 3, 4, 5, 9, 4, 4, 2, 3, 3, 2, 6, 3, 5, 3, 4, 3, 2, 2, 7, 1, 4, 8, 7, 4, 5, 3, 4, 3, 2, 5, 1, 3, 3, 2, 8, 3, 4, 2, 2, 6, 2, 2, 3, 4, 4, 4, 4, 2, 2, 6, 4, 5, 3, 4, 1, 2, 4, 2, 8, 3, 6, 5, 1, 3, 3, 2, 4, 2, 7, 9, 2, 4, 3, 2, 1, 1, 6, 7, 6, 3, 8, 8, 3, 2, 4, 6, 4, 1, 2, 2, 2, 2, 2, 3 };
        @(posedge clk);
        val = '{ 3, 5, 4, 3, 4, 5, 3, 4, 3, 4, 2, 5, 1, 2, 2, 6, 1, 3, 5, 2, 1, 3, 2, 4, 3, 2, 8, 1, 8, 2, 2, 3, 3, 2, 1, 3, 4, 3, 2, 9, 3, 9, 5, 4, 7, 1, 6, 2, 1, 1, 2, 3, 4, 3, 3, 1, 2, 1, 2, 3, 3, 3, 1, 6, 1, 2, 4, 3, 5, 5, 5, 2, 2, 7, 9, 5, 1, 2, 2, 8, 4, 3, 2, 4, 5, 3, 4, 5, 3, 3, 4, 3, 4, 2, 5, 7, 7, 4, 3, 2, 7, 2, 5, 3, 1, 4, 6, 2, 6, 6, 4, 3, 3, 4, 3, 2, 6, 4, 4, 5, 4, 2, 4, 1, 3, 2, 6, 5, 7, 6, 2, 1, 5, 4, 4, 8, 3, 4, 3, 6, 6, 3, 2, 4, 5, 1, 1, 2, 3, 3, 2, 3, 2, 4, 6, 3, 2, 3, 2, 4, 4, 1, 2, 1, 6, 3, 3, 5, 2, 6, 8, 2, 4, 6, 6, 8, 4, 5, 3, 3, 1, 2, 2, 2, 2, 2, 4, 6, 3, 2, 3, 6, 2, 3, 2, 4, 6, 3, 3, 3 };
        @(posedge clk);
        val = '{ 2, 4, 8, 5, 3, 8, 6, 6, 7, 4, 5, 5, 2, 4, 5, 4, 3, 1, 6, 2, 3, 3, 4, 2, 3, 7, 2, 7, 4, 2, 1, 4, 1, 2, 4, 4, 1, 1, 5, 1, 2, 6, 3, 4, 3, 3, 6, 3, 2, 2, 9, 2, 1, 3, 3, 2, 1, 3, 2, 3, 5, 4, 5, 7, 3, 2, 7, 4, 5, 5, 6, 1, 2, 5, 5, 5, 6, 2, 2, 2, 4, 4, 1, 6, 2, 2, 3, 5, 3, 2, 7, 3, 3, 4, 3, 2, 2, 4, 1, 2, 1, 4, 5, 8, 3, 5, 6, 2, 3, 3, 3, 5, 2, 4, 3, 5, 5, 4, 5, 2, 3, 2, 7, 2, 5, 1, 6, 3, 6, 5, 3, 3, 4, 6, 3, 3, 2, 7, 3, 3, 3, 3, 5, 4, 5, 6, 1, 2, 3, 2, 2, 5, 5, 2, 2, 2, 2, 6, 2, 8, 2, 2, 3, 4, 2, 3, 1, 6, 2, 4, 3, 3, 4, 2, 5, 7, 2, 3, 2, 2, 3, 1, 5, 2, 3, 2, 2, 8, 3, 2, 6, 5, 2, 2, 2, 6, 3, 4, 2, 2 };
        @(posedge clk);
        val = '{ 2, 2, 3, 3, 3, 1, 3, 6, 5, 4, 3, 3, 2, 6, 3, 2, 2, 1, 4, 2, 3, 3, 4, 2, 2, 2, 3, 4, 4, 2, 3, 4, 2, 3, 1, 2, 2, 2, 5, 5, 1, 6, 7, 4, 2, 2, 3, 1, 2, 2, 5, 2, 6, 4, 5, 3, 2, 2, 2, 5, 4, 2, 2, 3, 4, 2, 3, 7, 2, 3, 6, 4, 2, 2, 4, 6, 1, 2, 3, 4, 2, 1, 3, 5, 5, 1, 6, 6, 3, 3, 6, 2, 2, 3, 3, 2, 7, 5, 5, 2, 2, 8, 3, 4, 2, 7, 4, 6, 2, 6, 1, 5, 4, 2, 2, 1, 5, 7, 6, 3, 2, 4, 2, 2, 4, 2, 5, 5, 4, 5, 3, 2, 2, 5, 3, 3, 2, 5, 4, 4, 5, 3, 2, 6, 3, 3, 2, 2, 3, 2, 3, 2, 4, 3, 7, 6, 2, 2, 2, 3, 3, 1, 4, 2, 7, 2, 4, 6, 2, 3, 4, 4, 4, 6, 1, 7, 2, 3, 2, 2, 4, 1, 4, 3, 7, 2, 2, 5, 2, 3, 3, 4, 2, 2, 3, 2, 2, 4, 3, 4 };
        @(posedge clk);
        val = '{ 5, 4, 4, 4, 2, 3, 3, 4, 6, 3, 2, 6, 2, 3, 2, 3, 3, 2, 5, 2, 2, 1, 3, 2, 2, 8, 3, 1, 4, 5, 2, 4, 2, 2, 1, 5, 3, 7, 1, 8, 2, 7, 3, 5, 2, 3, 3, 3, 5, 2, 4, 3, 5, 3, 3, 2, 3, 2, 2, 4, 4, 3, 2, 2, 3, 2, 9, 8, 4, 3, 8, 4, 2, 5, 5, 8, 3, 5, 3, 5, 4, 2, 2, 7, 5, 5, 6, 3, 3, 3, 4, 3, 6, 4, 2, 6, 2, 4, 2, 2, 2, 5, 2, 3, 3, 3, 5, 5, 2, 2, 4, 3, 2, 4, 2, 1, 4, 2, 3, 5, 4, 3, 5, 1, 4, 2, 6, 3, 7, 2, 7, 5, 4, 6, 3, 5, 2, 7, 4, 1, 3, 3, 3, 3, 4, 2, 2, 2, 6, 2, 4, 5, 6, 2, 3, 3, 2, 2, 7, 4, 1, 1, 4, 2, 2, 2, 5, 6, 7, 2, 6, 4, 4, 5, 8, 9, 2, 3, 3, 1, 2, 2, 3, 6, 9, 2, 1, 1, 2, 4, 4, 3, 3, 1, 2, 3, 2, 4, 1, 2 };
        @(posedge clk);
        val = '{ 2, 5, 3, 4, 5, 4, 3, 2, 5, 2, 3, 7, 1, 4, 5, 2, 3, 2, 4, 2, 2, 2, 2, 2, 2, 3, 7, 3, 9, 2, 2, 4, 2, 2, 2, 5, 5, 2, 2, 2, 5, 5, 4, 2, 6, 5, 5, 4, 2, 2, 6, 3, 5, 2, 3, 2, 3, 4, 7, 3, 4, 2, 4, 5, 2, 1, 7, 2, 3, 8, 7, 4, 2, 6, 7, 8, 3, 2, 3, 2, 4, 2, 1, 6, 6, 3, 7, 4, 3, 2, 8, 7, 4, 3, 3, 7, 4, 5, 3, 2, 3, 5, 2, 2, 3, 4, 5, 2, 5, 5, 2, 2, 2, 1, 2, 3, 4, 4, 5, 4, 5, 2, 7, 2, 4, 4, 6, 4, 6, 3, 4, 2, 6, 2, 4, 3, 1, 3, 1, 6, 3, 3, 2, 2, 3, 1, 1, 2, 2, 4, 6, 3, 4, 2, 2, 2, 2, 4, 3, 1, 2, 2, 3, 2, 7, 3, 3, 3, 3, 6, 4, 7, 8, 5, 5, 4, 2, 4, 2, 2, 5, 3, 1, 4, 3, 2, 2, 3, 2, 2, 4, 4, 2, 1, 1, 4, 3, 2, 2, 6 };
        @(posedge clk);
        val = '{ 8, 4, 4, 3, 1, 2, 3, 2, 7, 5, 5, 2, 2, 7, 7, 2, 3, 1, 3, 2, 2, 2, 7, 4, 3, 4, 2, 3, 3, 2, 2, 3, 4, 3, 1, 3, 1, 2, 3, 8, 1, 6, 4, 3, 3, 2, 4, 2, 4, 3, 7, 1, 4, 1, 5, 1, 1, 1, 2, 4, 5, 4, 5, 4, 2, 3, 6, 9, 4, 2, 3, 2, 2, 2, 4, 7, 3, 1, 2, 4, 4, 2, 3, 5, 4, 7, 4, 3, 2, 2, 2, 5, 3, 2, 4, 1, 3, 2, 1, 2, 2, 5, 3, 4, 2, 4, 4, 3, 3, 5, 1, 3, 3, 2, 2, 6, 4, 4, 3, 1, 6, 2, 1, 2, 4, 2, 5, 7, 6, 4, 3, 2, 2, 2, 3, 3, 2, 4, 2, 2, 3, 3, 5, 4, 2, 3, 2, 1, 2, 4, 4, 6, 3, 3, 4, 4, 2, 3, 1, 5, 2, 2, 4, 2, 5, 3, 3, 6, 3, 6, 3, 2, 3, 4, 6, 8, 1, 2, 2, 2, 2, 2, 2, 2, 3, 2, 3, 3, 2, 3, 3, 1, 3, 2, 2, 4, 2, 2, 2, 2 };
        @(posedge clk);
        val = '{ 1, 4, 4, 3, 3, 2, 3, 6, 6, 4, 4, 3, 2, 6, 6, 3, 3, 2, 6, 2, 2, 3, 4, 3, 3, 3, 7, 3, 8, 2, 2, 4, 2, 3, 2, 3, 2, 1, 3, 5, 2, 5, 3, 2, 4, 7, 4, 2, 5, 1, 2, 2, 1, 5, 3, 2, 7, 3, 2, 4, 3, 2, 2, 9, 2, 2, 8, 3, 6, 4, 7, 2, 3, 5, 2, 4, 3, 3, 4, 6, 3, 1, 2, 3, 5, 2, 1, 5, 5, 4, 1, 4, 2, 5, 6, 2, 2, 5, 2, 1, 2, 5, 2, 4, 3, 4, 5, 2, 5, 5, 4, 4, 2, 4, 3, 6, 5, 5, 5, 2, 2, 3, 4, 2, 3, 2, 6, 7, 5, 4, 4, 3, 2, 5, 4, 3, 2, 5, 5, 2, 3, 3, 1, 2, 4, 2, 2, 1, 3, 2, 1, 2, 3, 4, 4, 5, 3, 2, 4, 5, 2, 1, 4, 3, 8, 3, 3, 5, 2, 4, 2, 2, 3, 6, 7, 4, 3, 1, 5, 2, 2, 2, 1, 3, 5, 2, 2, 2, 4, 2, 5, 3, 2, 3, 2, 2, 4, 3, 3, 5 };
        @(posedge clk);
        val = '{ 5, 2, 2, 6, 2, 4, 6, 7, 8, 3, 4, 1, 2, 1, 2, 3, 3, 2, 4, 3, 2, 2, 3, 5, 3, 2, 2, 3, 4, 2, 2, 4, 2, 3, 2, 4, 2, 4, 3, 5, 2, 4, 3, 7, 6, 2, 3, 3, 3, 2, 4, 2, 4, 2, 6, 2, 1, 2, 3, 4, 4, 1, 2, 3, 4, 4, 9, 4, 2, 3, 1, 3, 1, 4, 2, 4, 3, 2, 5, 2, 3, 2, 2, 5, 3, 3, 1, 2, 2, 3, 6, 3, 3, 4, 2, 2, 2, 4, 1, 1, 3, 2, 3, 4, 7, 4, 5, 2, 5, 9, 3, 3, 2, 1, 3, 4, 4, 4, 5, 1, 4, 3, 3, 3, 1, 4, 1, 6, 4, 2, 4, 6, 4, 2, 2, 3, 3, 4, 2, 7, 2, 2, 3, 5, 4, 3, 1, 1, 3, 2, 4, 5, 5, 2, 6, 7, 3, 3, 6, 2, 2, 2, 4, 1, 5, 3, 6, 4, 2, 1, 5, 4, 3, 5, 3, 3, 4, 6, 1, 2, 2, 2, 5, 7, 6, 2, 2, 3, 2, 3, 4, 4, 3, 1, 1, 5, 3, 2, 4, 2 };
        @(posedge clk);
        val = '{ 6, 7, 4, 2, 4, 4, 3, 1, 3, 3, 5, 5, 2, 2, 3, 3, 6, 4, 3, 2, 3, 3, 5, 2, 1, 5, 3, 2, 6, 2, 2, 4, 2, 3, 2, 4, 6, 2, 3, 5, 1, 5, 6, 3, 4, 2, 3, 4, 2, 4, 6, 2, 3, 3, 3, 2, 6, 2, 2, 4, 4, 5, 1, 3, 2, 2, 5, 2, 4, 3, 4, 1, 3, 2, 2, 8, 8, 2, 1, 2, 5, 2, 1, 5, 3, 1, 3, 2, 3, 3, 8, 2, 3, 2, 5, 8, 2, 5, 2, 1, 2, 5, 2, 2, 3, 5, 6, 2, 2, 2, 4, 3, 1, 2, 3, 2, 5, 2, 6, 2, 3, 2, 2, 2, 1, 4, 6, 6, 4, 2, 2, 2, 2, 6, 3, 3, 2, 5, 4, 5, 4, 3, 4, 6, 1, 2, 4, 3, 2, 2, 4, 7, 3, 4, 1, 3, 4, 2, 4, 4, 1, 1, 3, 2, 2, 2, 2, 8, 3, 2, 3, 2, 4, 2, 3, 8, 6, 4, 2, 2, 2, 3, 3, 3, 1, 2, 2, 4, 3, 3, 1, 2, 2, 2, 2, 6, 6, 7, 3, 5 };
        @(posedge clk);
        val = '{ 2, 5, 6, 3, 6, 1, 6, 6, 9, 3, 4, 5, 2, 2, 8, 3, 3, 2, 5, 4, 3, 3, 4, 3, 1, 2, 4, 2, 7, 1, 2, 3, 4, 3, 1, 4, 7, 4, 3, 4, 2, 6, 6, 1, 2, 3, 2, 3, 5, 2, 3, 5, 3, 3, 1, 2, 5, 9, 1, 7, 4, 3, 3, 7, 5, 3, 1, 3, 5, 7, 1, 1, 2, 9, 4, 7, 2, 2, 4, 4, 1, 4, 2, 8, 2, 3, 2, 4, 3, 3, 2, 5, 4, 3, 4, 2, 2, 9, 2, 2, 2, 8, 3, 4, 3, 4, 2, 2, 2, 2, 2, 5, 2, 2, 5, 4, 1, 6, 4, 4, 3, 1, 7, 2, 6, 2, 5, 9, 5, 5, 6, 4, 5, 5, 2, 3, 4, 4, 2, 6, 5, 4, 1, 4, 3, 2, 2, 1, 3, 2, 4, 2, 3, 2, 4, 6, 4, 3, 3, 1, 2, 2, 4, 3, 8, 3, 5, 4, 2, 2, 1, 1, 5, 6, 3, 9, 3, 4, 2, 2, 2, 2, 3, 3, 6, 2, 3, 9, 3, 2, 5, 4, 2, 2, 2, 4, 2, 2, 3, 4 };
        @(posedge clk);
        val = '{ 2, 2, 1, 6, 1, 3, 3, 2, 8, 3, 2, 5, 3, 3, 4, 2, 3, 2, 3, 3, 3, 3, 3, 2, 2, 5, 3, 8, 4, 3, 1, 4, 2, 3, 4, 7, 6, 2, 3, 4, 3, 6, 2, 5, 4, 1, 2, 3, 3, 1, 6, 2, 4, 4, 3, 1, 2, 1, 2, 5, 2, 3, 4, 5, 2, 2, 3, 7, 2, 4, 3, 2, 2, 7, 2, 6, 3, 4, 3, 3, 2, 1, 2, 9, 4, 2, 1, 3, 3, 3, 6, 6, 2, 3, 3, 3, 1, 2, 1, 1, 3, 4, 3, 6, 3, 2, 6, 2, 3, 8, 3, 3, 2, 4, 2, 2, 5, 4, 6, 2, 1, 3, 4, 2, 3, 3, 3, 5, 8, 5, 3, 2, 1, 5, 3, 5, 2, 4, 3, 2, 4, 3, 2, 3, 4, 3, 2, 1, 2, 2, 2, 6, 4, 1, 7, 3, 4, 6, 2, 2, 2, 2, 5, 3, 4, 3, 5, 5, 3, 3, 2, 2, 4, 8, 2, 6, 1, 3, 1, 4, 5, 2, 2, 3, 4, 2, 2, 3, 2, 2, 4, 4, 2, 2, 2, 6, 2, 3, 4, 2 };
        @(posedge clk);
        val = '{ 4, 4, 3, 4, 5, 7, 3, 2, 5, 4, 3, 2, 2, 5, 5, 3, 2, 2, 5, 2, 3, 4, 3, 4, 1, 4, 3, 2, 5, 3, 1, 3, 2, 2, 3, 4, 2, 5, 2, 7, 3, 6, 4, 6, 2, 2, 6, 2, 4, 2, 4, 2, 2, 2, 3, 2, 3, 1, 1, 2, 2, 2, 4, 8, 3, 1, 5, 2, 2, 4, 2, 3, 3, 4, 4, 6, 4, 2, 2, 2, 6, 2, 2, 6, 5, 4, 7, 5, 2, 3, 2, 7, 4, 3, 2, 6, 2, 5, 3, 2, 2, 5, 5, 6, 3, 4, 6, 2, 3, 5, 3, 2, 4, 2, 3, 7, 5, 1, 5, 5, 3, 3, 3, 2, 2, 1, 5, 6, 4, 4, 4, 2, 2, 3, 2, 3, 2, 3, 3, 1, 2, 4, 2, 6, 2, 5, 2, 3, 5, 1, 4, 4, 3, 1, 6, 4, 2, 6, 2, 2, 1, 1, 4, 2, 4, 3, 5, 5, 2, 3, 4, 4, 5, 4, 6, 5, 2, 1, 1, 4, 2, 2, 7, 2, 8, 2, 4, 2, 3, 3, 6, 5, 2, 1, 2, 7, 3, 6, 3, 4 };
        @(posedge clk);
        val = '{ 1, 2, 7, 2, 3, 5, 3, 2, 5, 2, 5, 2, 2, 4, 3, 3, 1, 2, 5, 2, 2, 5, 2, 2, 3, 8, 3, 4, 4, 2, 2, 4, 2, 2, 4, 5, 2, 2, 2, 5, 3, 6, 3, 1, 2, 2, 6, 2, 2, 2, 3, 2, 7, 2, 2, 1, 2, 1, 7, 3, 3, 3, 1, 6, 1, 2, 6, 3, 3, 5, 6, 2, 1, 8, 2, 2, 3, 2, 3, 8, 3, 2, 2, 7, 5, 3, 6, 6, 2, 4, 4, 5, 3, 3, 2, 9, 4, 2, 2, 2, 8, 5, 5, 3, 5, 4, 6, 4, 5, 9, 3, 3, 1, 2, 2, 2, 2, 4, 6, 2, 3, 3, 2, 2, 5, 1, 6, 8, 4, 3, 5, 2, 3, 4, 3, 3, 2, 3, 1, 3, 4, 3, 2, 2, 4, 4, 1, 2, 2, 2, 3, 4, 4, 5, 4, 3, 4, 1, 2, 3, 2, 2, 4, 2, 2, 8, 1, 7, 2, 3, 1, 2, 5, 2, 6, 6, 1, 3, 1, 2, 2, 1, 2, 3, 6, 2, 1, 4, 1, 3, 5, 3, 1, 1, 2, 6, 2, 3, 3, 3 };
        @(posedge clk);
        val = '{ 3, 4, 5, 3, 3, 4, 3, 2, 6, 2, 3, 2, 5, 2, 2, 1, 3, 2, 8, 2, 2, 2, 3, 2, 3, 2, 6, 2, 7, 2, 2, 4, 1, 5, 2, 3, 7, 4, 4, 5, 2, 5, 4, 7, 2, 4, 2, 4, 8, 4, 3, 1, 7, 3, 3, 2, 2, 2, 4, 4, 2, 2, 2, 3, 1, 2, 6, 2, 2, 3, 4, 1, 2, 5, 5, 5, 3, 3, 4, 3, 6, 2, 2, 8, 5, 2, 5, 4, 3, 2, 5, 6, 3, 5, 1, 2, 4, 3, 4, 1, 5, 5, 3, 3, 4, 3, 7, 3, 2, 2, 3, 3, 3, 3, 3, 2, 6, 4, 4, 3, 9, 1, 3, 2, 5, 3, 6, 6, 2, 5, 5, 2, 2, 2, 3, 3, 2, 5, 7, 2, 6, 3, 2, 3, 4, 2, 2, 2, 1, 4, 2, 5, 3, 3, 1, 1, 4, 4, 2, 4, 2, 2, 2, 3, 2, 3, 6, 3, 2, 3, 3, 1, 4, 1, 4, 9, 6, 4, 3, 3, 4, 3, 2, 6, 5, 2, 1, 5, 1, 3, 3, 2, 2, 3, 2, 7, 2, 5, 2, 4 };
        @(posedge clk);
        val = '{ 2, 4, 6, 3, 5, 5, 5, 4, 7, 3, 4, 5, 3, 2, 3, 3, 3, 3, 9, 1, 2, 4, 1, 2, 3, 4, 5, 4, 5, 1, 2, 3, 3, 1, 3, 6, 2, 3, 3, 7, 2, 9, 4, 2, 4, 2, 4, 5, 3, 3, 3, 2, 6, 7, 2, 2, 1, 2, 3, 5, 4, 1, 3, 7, 3, 1, 2, 5, 3, 3, 7, 1, 2, 4, 3, 5, 2, 2, 2, 1, 2, 3, 2, 5, 5, 2, 1, 5, 3, 1, 4, 2, 1, 2, 4, 4, 3, 5, 2, 3, 2, 6, 2, 4, 6, 5, 6, 3, 3, 9, 3, 3, 2, 2, 3, 7, 4, 4, 3, 3, 4, 2, 7, 2, 5, 2, 4, 6, 8, 4, 2, 3, 4, 5, 3, 3, 1, 4, 2, 1, 3, 3, 7, 6, 1, 4, 1, 2, 5, 3, 4, 6, 6, 6, 5, 5, 3, 4, 2, 2, 2, 1, 4, 3, 2, 4, 5, 5, 1, 4, 2, 2, 3, 3, 3, 6, 1, 4, 4, 2, 5, 2, 4, 3, 5, 2, 2, 3, 2, 2, 4, 3, 2, 2, 2, 7, 3, 3, 2, 3 };
        @(posedge clk);
        val = '{ 2, 3, 2, 3, 3, 4, 3, 2, 9, 1, 4, 2, 2, 3, 4, 3, 4, 4, 7, 2, 1, 5, 5, 1, 3, 3, 2, 7, 4, 3, 3, 4, 2, 5, 2, 2, 2, 2, 4, 4, 4, 4, 4, 2, 5, 7, 2, 5, 2, 2, 6, 3, 5, 2, 4, 2, 2, 2, 4, 5, 4, 3, 3, 4, 2, 4, 5, 8, 4, 6, 7, 2, 2, 6, 5, 6, 9, 2, 2, 2, 3, 4, 1, 7, 4, 2, 4, 3, 1, 3, 4, 3, 4, 4, 4, 5, 2, 4, 3, 5, 5, 8, 2, 5, 4, 5, 6, 4, 3, 5, 3, 3, 3, 3, 3, 5, 6, 4, 5, 4, 3, 2, 4, 2, 2, 3, 6, 5, 5, 5, 5, 2, 3, 6, 4, 3, 1, 4, 3, 2, 7, 4, 4, 2, 1, 2, 1, 2, 3, 2, 3, 4, 1, 3, 7, 6, 4, 6, 2, 6, 2, 3, 4, 3, 6, 2, 3, 5, 2, 5, 7, 1, 3, 7, 4, 8, 4, 7, 2, 2, 2, 2, 1, 2, 4, 2, 4, 4, 2, 3, 4, 4, 2, 1, 2, 3, 9, 3, 3, 3 };
        @(posedge clk);
        val = '{ 4, 4, 2, 3, 4, 5, 4, 2, 5, 3, 5, 2, 2, 3, 4, 3, 2, 4, 3, 2, 3, 5, 3, 2, 4, 4, 1, 9, 4, 2, 2, 2, 2, 2, 2, 6, 2, 4, 5, 3, 3, 6, 2, 5, 3, 2, 2, 1, 2, 2, 4, 4, 6, 5, 3, 3, 2, 2, 8, 2, 4, 3, 2, 6, 3, 2, 2, 5, 4, 3, 3, 3, 1, 8, 6, 3, 3, 3, 2, 3, 5, 1, 2, 8, 5, 2, 3, 5, 3, 2, 2, 2, 1, 3, 6, 4, 3, 5, 2, 2, 1, 5, 2, 2, 2, 3, 6, 2, 3, 7, 2, 3, 2, 3, 3, 6, 4, 1, 3, 2, 5, 3, 2, 1, 5, 2, 1, 4, 5, 4, 4, 5, 5, 5, 1, 3, 2, 3, 4, 3, 2, 3, 2, 3, 4, 3, 4, 1, 3, 7, 4, 4, 3, 2, 1, 3, 7, 2, 5, 3, 2, 2, 2, 4, 4, 3, 3, 2, 2, 3, 2, 2, 5, 7, 4, 5, 4, 1, 2, 3, 4, 1, 2, 2, 4, 2, 2, 3, 3, 2, 5, 2, 1, 2, 1, 5, 2, 3, 2, 3 };
        @(posedge clk);
        val = '{ 3, 6, 3, 3, 2, 1, 1, 2, 4, 3, 4, 3, 1, 7, 3, 3, 1, 1, 7, 2, 3, 4, 3, 1, 3, 3, 2, 2, 5, 2, 2, 4, 2, 3, 2, 2, 6, 1, 5, 4, 2, 5, 6, 1, 6, 2, 3, 4, 5, 2, 4, 2, 5, 2, 4, 1, 2, 1, 2, 5, 2, 5, 5, 3, 2, 2, 3, 8, 1, 3, 8, 2, 4, 4, 7, 4, 5, 2, 4, 2, 2, 2, 2, 8, 8, 2, 5, 3, 2, 3, 2, 3, 1, 2, 5, 3, 2, 2, 2, 2, 5, 6, 3, 4, 3, 3, 5, 2, 3, 4, 3, 3, 1, 2, 3, 5, 5, 6, 3, 5, 4, 1, 6, 2, 4, 3, 6, 4, 8, 2, 3, 4, 3, 6, 4, 2, 4, 4, 3, 3, 3, 4, 6, 4, 4, 2, 2, 8, 2, 2, 3, 4, 3, 4, 6, 2, 7, 5, 3, 3, 3, 3, 1, 2, 5, 3, 3, 3, 3, 5, 2, 2, 4, 2, 4, 7, 2, 4, 2, 2, 4, 3, 2, 3, 2, 2, 2, 9, 3, 3, 4, 4, 2, 2, 1, 6, 2, 3, 5, 8 };
        @(posedge clk);
        val = '{ 4, 5, 3, 1, 3, 6, 3, 5, 7, 2, 3, 4, 2, 2, 1, 3, 3, 5, 4, 2, 1, 5, 4, 5, 3, 1, 4, 3, 3, 3, 2, 3, 2, 2, 1, 4, 3, 2, 3, 7, 2, 4, 3, 5, 2, 3, 6, 6, 3, 3, 8, 3, 5, 4, 3, 2, 3, 2, 2, 2, 2, 4, 1, 4, 3, 2, 3, 5, 2, 4, 6, 2, 2, 5, 9, 3, 3, 3, 4, 3, 2, 2, 3, 7, 5, 4, 1, 6, 3, 3, 2, 6, 2, 2, 2, 4, 5, 4, 6, 2, 2, 5, 4, 3, 2, 2, 5, 5, 5, 4, 2, 3, 2, 3, 3, 3, 5, 4, 5, 3, 5, 1, 3, 2, 4, 1, 3, 4, 4, 5, 4, 3, 5, 3, 4, 4, 2, 5, 2, 4, 8, 1, 2, 3, 2, 2, 3, 2, 8, 1, 4, 6, 1, 3, 7, 3, 3, 5, 1, 5, 3, 3, 2, 1, 6, 1, 2, 6, 5, 4, 2, 1, 3, 6, 8, 8, 2, 3, 2, 1, 1, 2, 3, 6, 6, 2, 1, 3, 3, 3, 3, 4, 2, 3, 2, 2, 4, 6, 1, 5 };
        @(posedge clk);
        val = '{ 8, 1, 3, 5, 1, 4, 2, 4, 5, 4, 4, 5, 1, 1, 7, 1, 3, 2, 4, 2, 2, 3, 3, 4, 3, 3, 3, 9, 5, 2, 2, 4, 1, 1, 2, 4, 5, 2, 2, 4, 2, 4, 5, 4, 4, 3, 3, 2, 3, 2, 4, 3, 4, 2, 2, 2, 2, 2, 2, 2, 4, 2, 2, 5, 4, 2, 3, 3, 3, 4, 3, 4, 2, 5, 2, 3, 3, 2, 2, 3, 3, 2, 2, 8, 6, 4, 6, 3, 2, 3, 2, 2, 4, 3, 3, 8, 2, 5, 2, 2, 8, 5, 4, 5, 2, 4, 5, 2, 2, 4, 6, 3, 4, 2, 3, 2, 3, 4, 5, 2, 6, 2, 4, 2, 5, 5, 4, 2, 5, 4, 6, 2, 5, 3, 2, 2, 4, 2, 4, 3, 5, 3, 2, 3, 3, 2, 2, 2, 5, 2, 2, 4, 6, 4, 7, 3, 2, 5, 3, 2, 2, 2, 2, 2, 6, 3, 2, 4, 2, 3, 2, 6, 9, 9, 7, 6, 2, 6, 2, 2, 5, 3, 4, 8, 2, 2, 3, 8, 4, 3, 4, 2, 3, 7, 2, 3, 7, 6, 5, 2 };
        @(posedge clk);
        val = '{ 4, 5, 8, 1, 3, 6, 3, 3, 6, 4, 3, 4, 2, 5, 7, 3, 3, 2, 7, 2, 4, 8, 4, 3, 2, 7, 1, 5, 6, 3, 2, 4, 4, 2, 1, 3, 1, 2, 3, 7, 1, 2, 2, 2, 7, 2, 3, 3, 2, 2, 2, 2, 4, 4, 4, 2, 7, 1, 4, 5, 4, 2, 5, 4, 3, 3, 7, 6, 5, 3, 5, 2, 3, 7, 4, 8, 4, 2, 4, 3, 3, 2, 2, 5, 6, 3, 7, 3, 3, 3, 6, 5, 4, 3, 2, 5, 3, 3, 3, 2, 7, 5, 1, 3, 6, 4, 5, 3, 5, 8, 3, 3, 1, 2, 3, 6, 2, 4, 2, 4, 3, 2, 4, 6, 7, 1, 5, 9, 7, 2, 4, 2, 3, 2, 3, 3, 5, 5, 2, 4, 5, 2, 2, 4, 3, 7, 2, 2, 3, 2, 4, 3, 4, 2, 7, 9, 2, 3, 1, 8, 2, 1, 4, 2, 8, 3, 3, 6, 1, 8, 3, 1, 2, 6, 6, 9, 2, 4, 4, 1, 3, 2, 3, 7, 2, 2, 2, 3, 2, 3, 3, 2, 1, 2, 3, 2, 5, 2, 4, 3 };
        @(posedge clk);
        val = '{ 8, 6, 7, 2, 2, 5, 3, 5, 4, 1, 5, 3, 2, 4, 2, 5, 4, 3, 5, 1, 3, 2, 3, 2, 3, 4, 7, 4, 5, 2, 2, 3, 4, 3, 6, 3, 2, 2, 5, 5, 1, 5, 5, 6, 4, 4, 2, 5, 7, 2, 4, 3, 4, 3, 2, 2, 2, 2, 2, 3, 4, 8, 2, 4, 2, 1, 4, 4, 6, 3, 3, 4, 1, 4, 3, 5, 7, 2, 1, 5, 4, 4, 3, 5, 5, 3, 1, 3, 4, 5, 3, 3, 4, 2, 5, 7, 6, 4, 2, 3, 6, 3, 4, 2, 4, 2, 5, 2, 5, 7, 2, 3, 2, 2, 3, 2, 3, 4, 6, 1, 4, 4, 5, 2, 2, 2, 3, 5, 3, 5, 7, 3, 2, 4, 4, 3, 1, 5, 4, 5, 2, 4, 2, 5, 1, 2, 3, 3, 2, 3, 5, 5, 4, 2, 5, 2, 3, 6, 4, 6, 2, 3, 2, 2, 4, 2, 3, 5, 3, 5, 8, 2, 7, 6, 8, 8, 4, 4, 2, 2, 2, 2, 4, 5, 3, 2, 3, 6, 3, 3, 5, 3, 2, 3, 4, 5, 4, 1, 2, 1 };
        @(posedge clk);
        val = '{ 3, 4, 2, 2, 2, 3, 3, 3, 2, 2, 3, 5, 2, 2, 2, 3, 2, 3, 4, 2, 1, 5, 1, 2, 2, 8, 3, 5, 5, 2, 2, 2, 3, 3, 2, 3, 2, 1, 1, 4, 7, 7, 3, 7, 3, 2, 2, 5, 5, 2, 5, 3, 4, 2, 6, 2, 2, 2, 2, 3, 3, 4, 4, 8, 3, 6, 6, 4, 2, 3, 8, 2, 2, 8, 6, 9, 4, 1, 3, 3, 4, 2, 2, 8, 6, 2, 6, 4, 2, 2, 8, 2, 4, 2, 1, 6, 2, 7, 1, 2, 4, 1, 1, 5, 3, 4, 7, 3, 3, 3, 3, 3, 2, 3, 3, 2, 4, 4, 7, 5, 3, 2, 6, 2, 3, 3, 5, 9, 5, 3, 5, 7, 4, 1, 3, 4, 2, 4, 4, 3, 4, 7, 1, 6, 2, 2, 3, 2, 3, 2, 6, 6, 2, 5, 2, 6, 3, 3, 7, 1, 1, 1, 5, 1, 7, 3, 5, 5, 2, 3, 3, 3, 3, 6, 3, 8, 2, 2, 2, 2, 3, 1, 4, 9, 3, 1, 2, 2, 2, 3, 4, 4, 2, 2, 2, 5, 1, 3, 7, 3 };
        @(posedge clk);
        val = '{ 2, 4, 2, 3, 2, 5, 3, 1, 5, 1, 4, 8, 1, 2, 7, 5, 5, 2, 8, 2, 2, 3, 5, 1, 2, 2, 3, 4, 5, 2, 1, 3, 2, 2, 2, 4, 2, 2, 4, 6, 3, 4, 4, 7, 4, 5, 1, 3, 4, 2, 4, 2, 5, 3, 4, 2, 3, 2, 2, 2, 5, 4, 4, 9, 5, 6, 9, 9, 2, 4, 2, 1, 7, 6, 3, 3, 3, 2, 4, 3, 4, 2, 1, 8, 5, 7, 6, 5, 4, 3, 7, 3, 4, 3, 2, 2, 2, 9, 5, 2, 3, 5, 8, 3, 3, 4, 7, 4, 3, 5, 8, 3, 3, 3, 2, 6, 5, 3, 3, 3, 4, 3, 4, 2, 6, 2, 4, 5, 7, 2, 3, 6, 2, 3, 2, 3, 2, 5, 4, 2, 6, 2, 4, 6, 2, 2, 2, 2, 2, 2, 3, 1, 3, 2, 8, 4, 1, 4, 2, 2, 3, 1, 2, 3, 7, 2, 5, 9, 2, 5, 2, 4, 5, 6, 4, 5, 4, 4, 2, 2, 2, 3, 2, 6, 3, 2, 1, 3, 5, 3, 4, 4, 1, 1, 2, 6, 2, 5, 4, 3 };
        @(posedge clk);
        val = '{ 3, 4, 3, 2, 3, 6, 4, 6, 5, 6, 2, 4, 3, 2, 6, 3, 3, 1, 6, 2, 2, 2, 3, 2, 2, 5, 2, 1, 6, 2, 3, 2, 3, 1, 2, 4, 2, 5, 4, 6, 4, 4, 6, 2, 4, 2, 3, 5, 2, 1, 4, 3, 4, 2, 3, 2, 2, 1, 3, 7, 4, 3, 5, 6, 3, 2, 3, 3, 2, 6, 6, 1, 3, 7, 3, 5, 3, 2, 3, 3, 6, 3, 1, 5, 2, 3, 7, 9, 3, 2, 2, 6, 4, 3, 2, 3, 4, 5, 4, 2, 1, 3, 4, 4, 5, 3, 3, 4, 4, 8, 4, 3, 2, 1, 3, 1, 5, 4, 6, 2, 1, 2, 3, 2, 2, 2, 6, 6, 9, 2, 4, 2, 4, 5, 2, 2, 2, 3, 4, 7, 9, 3, 2, 4, 2, 3, 2, 2, 8, 3, 3, 3, 2, 3, 1, 5, 3, 6, 7, 3, 2, 2, 4, 2, 4, 4, 8, 3, 2, 3, 4, 2, 4, 8, 4, 5, 2, 4, 4, 2, 3, 4, 2, 3, 2, 2, 2, 3, 3, 3, 3, 2, 2, 2, 8, 7, 3, 2, 4, 2 };
        @(posedge clk);
        val = '{ 3, 2, 2, 2, 3, 4, 5, 5, 2, 2, 4, 5, 2, 1, 2, 3, 3, 3, 7, 2, 5, 5, 1, 4, 3, 3, 7, 6, 9, 3, 3, 3, 3, 5, 2, 4, 3, 3, 3, 4, 2, 3, 4, 7, 4, 3, 5, 3, 5, 4, 7, 4, 7, 5, 3, 2, 2, 2, 2, 4, 6, 3, 2, 3, 2, 2, 2, 4, 2, 2, 5, 3, 2, 3, 5, 8, 3, 2, 2, 3, 3, 2, 2, 6, 3, 1, 7, 4, 3, 2, 2, 8, 5, 2, 5, 8, 6, 5, 2, 5, 2, 8, 3, 5, 3, 4, 6, 2, 2, 5, 8, 2, 3, 4, 4, 5, 2, 4, 4, 2, 1, 2, 3, 1, 6, 2, 5, 7, 7, 5, 4, 2, 4, 3, 3, 3, 4, 5, 1, 3, 5, 3, 2, 4, 2, 4, 2, 2, 3, 4, 4, 4, 3, 3, 3, 2, 3, 3, 3, 3, 2, 2, 3, 4, 6, 3, 2, 4, 2, 3, 3, 2, 4, 6, 6, 6, 2, 6, 3, 2, 5, 3, 4, 2, 3, 2, 1, 4, 5, 2, 4, 3, 3, 2, 2, 7, 3, 3, 4, 2 };
        @(posedge clk);
        val = '{ 4, 1, 4, 3, 4, 3, 5, 3, 3, 3, 5, 3, 2, 3, 3, 4, 3, 2, 3, 1, 1, 2, 3, 2, 4, 7, 6, 4, 4, 2, 2, 4, 2, 3, 1, 6, 4, 4, 5, 6, 5, 6, 4, 3, 2, 2, 5, 4, 3, 2, 2, 1, 5, 2, 3, 1, 2, 2, 2, 2, 5, 4, 4, 4, 2, 2, 6, 4, 2, 2, 8, 5, 2, 5, 3, 3, 3, 2, 4, 2, 2, 3, 4, 8, 4, 3, 2, 6, 3, 1, 2, 1, 2, 3, 3, 4, 5, 2, 2, 2, 4, 5, 3, 2, 4, 3, 5, 4, 4, 8, 3, 3, 2, 8, 6, 2, 6, 6, 5, 3, 2, 3, 5, 3, 4, 4, 4, 3, 8, 4, 4, 3, 2, 3, 3, 2, 2, 8, 3, 6, 7, 7, 1, 3, 2, 2, 2, 2, 6, 2, 3, 1, 7, 4, 2, 3, 3, 4, 4, 4, 2, 2, 1, 2, 7, 3, 3, 5, 2, 4, 4, 2, 5, 8, 7, 6, 2, 4, 2, 1, 4, 2, 2, 5, 4, 2, 2, 7, 2, 3, 4, 3, 3, 3, 2, 7, 2, 2, 7, 5 };
        @(posedge clk);
        val = '{ 2, 5, 2, 3, 3, 1, 4, 4, 7, 2, 3, 4, 2, 6, 2, 2, 5, 3, 6, 2, 3, 2, 4, 2, 4, 2, 3, 5, 4, 3, 1, 5, 4, 4, 2, 6, 1, 3, 4, 5, 2, 4, 2, 7, 4, 2, 6, 5, 5, 1, 5, 4, 3, 3, 3, 2, 4, 2, 3, 4, 1, 1, 6, 6, 2, 2, 4, 5, 2, 7, 2, 6, 2, 9, 5, 6, 4, 2, 2, 5, 2, 2, 2, 5, 7, 2, 5, 3, 2, 2, 6, 7, 6, 5, 5, 5, 7, 3, 1, 2, 4, 3, 2, 8, 3, 4, 5, 3, 5, 9, 3, 2, 5, 3, 3, 2, 3, 2, 7, 6, 5, 3, 2, 2, 7, 2, 5, 6, 7, 4, 4, 7, 2, 2, 2, 3, 4, 5, 4, 2, 3, 3, 1, 4, 2, 6, 2, 2, 2, 8, 2, 4, 3, 2, 6, 5, 5, 4, 2, 1, 3, 1, 3, 2, 5, 4, 2, 4, 2, 4, 3, 2, 9, 6, 3, 9, 5, 4, 3, 2, 6, 2, 2, 5, 8, 1, 6, 4, 2, 3, 2, 4, 3, 3, 2, 6, 1, 3, 2, 5 };
        @(posedge clk);
        val = '{ 8, 6, 8, 4, 3, 6, 4, 7, 6, 4, 6, 4, 2, 2, 5, 3, 2, 2, 2, 2, 1, 2, 2, 2, 3, 2, 3, 2, 4, 2, 2, 3, 2, 2, 2, 4, 6, 4, 4, 8, 2, 5, 3, 1, 4, 3, 5, 5, 8, 2, 6, 2, 3, 5, 6, 2, 1, 2, 2, 3, 5, 3, 7, 2, 3, 5, 8, 6, 4, 2, 6, 7, 2, 7, 3, 4, 3, 1, 3, 3, 4, 4, 2, 8, 6, 6, 7, 4, 3, 3, 4, 3, 4, 2, 3, 6, 2, 3, 2, 2, 2, 7, 3, 2, 3, 2, 5, 2, 2, 5, 4, 4, 2, 3, 3, 5, 2, 2, 4, 2, 3, 2, 3, 2, 6, 2, 6, 5, 3, 4, 7, 2, 2, 1, 4, 3, 4, 4, 2, 1, 2, 3, 2, 6, 5, 5, 1, 3, 9, 1, 2, 4, 2, 5, 2, 2, 1, 7, 2, 2, 3, 2, 3, 2, 2, 7, 3, 6, 2, 1, 4, 3, 7, 8, 3, 8, 1, 4, 3, 2, 3, 1, 3, 4, 7, 2, 2, 6, 3, 3, 3, 2, 2, 2, 2, 7, 3, 3, 2, 2 };
        @(posedge clk);
        val = '{ 5, 4, 5, 3, 2, 5, 2, 2, 5, 5, 4, 2, 4, 1, 3, 3, 2, 3, 9, 2, 2, 3, 2, 2, 4, 4, 3, 2, 3, 2, 2, 2, 1, 3, 3, 3, 2, 2, 1, 3, 2, 6, 6, 3, 5, 4, 5, 3, 2, 2, 5, 2, 4, 2, 3, 3, 2, 2, 3, 4, 1, 4, 8, 9, 3, 2, 4, 5, 2, 5, 2, 8, 1, 7, 2, 3, 5, 2, 2, 2, 2, 4, 1, 7, 4, 2, 8, 6, 4, 4, 4, 7, 2, 2, 7, 8, 4, 9, 7, 2, 8, 5, 1, 4, 4, 2, 3, 3, 4, 8, 2, 4, 5, 7, 3, 4, 2, 8, 5, 2, 2, 2, 4, 2, 4, 3, 6, 1, 6, 4, 3, 4, 1, 3, 1, 2, 2, 5, 2, 2, 1, 3, 4, 5, 3, 3, 1, 4, 5, 2, 3, 5, 4, 2, 2, 5, 5, 8, 2, 4, 2, 3, 2, 1, 2, 4, 3, 6, 3, 1, 2, 4, 3, 8, 3, 9, 2, 3, 2, 3, 2, 2, 2, 3, 2, 2, 2, 4, 2, 2, 5, 4, 4, 3, 1, 6, 5, 6, 2, 3 };
        @(posedge clk);
        val = '{ 2, 3, 3, 2, 1, 6, 4, 6, 7, 3, 4, 2, 2, 2, 6, 2, 2, 3, 9, 1, 5, 4, 2, 1, 1, 2, 3, 4, 4, 1, 2, 4, 3, 2, 3, 6, 1, 2, 4, 6, 4, 4, 5, 3, 4, 3, 6, 2, 4, 2, 7, 2, 5, 1, 3, 2, 2, 2, 2, 3, 3, 4, 9, 7, 2, 2, 3, 2, 4, 9, 2, 9, 3, 7, 5, 8, 2, 2, 3, 5, 4, 3, 1, 5, 2, 3, 9, 4, 1, 2, 4, 6, 3, 2, 1, 2, 2, 5, 3, 6, 6, 3, 2, 5, 6, 4, 5, 3, 4, 8, 2, 3, 2, 4, 2, 2, 4, 4, 2, 3, 3, 2, 3, 7, 5, 3, 7, 5, 3, 5, 3, 1, 4, 5, 5, 4, 3, 3, 2, 5, 3, 3, 3, 3, 3, 5, 2, 3, 2, 2, 4, 4, 5, 2, 9, 2, 2, 9, 2, 3, 2, 2, 4, 2, 4, 6, 3, 4, 2, 6, 6, 2, 3, 6, 5, 9, 2, 2, 2, 2, 1, 1, 3, 7, 7, 2, 5, 2, 4, 3, 3, 2, 2, 2, 2, 1, 3, 4, 4, 1 };
        @(posedge clk);

        // done storing
        bank_en = 0;
        val = '0;

        repeat (500) @(posedge clk);

        $finish;
    end

endmodule
