
`timescale 1ns/1ps

module tb_puzzle1;

    localparam MAX_LENGTH = 10;
    localparam SUM_SIZE   = 50;
    localparam NUM_RANGES = 30;

    logic clk;
    logic rst_n;
    logic vld;

    logic [NUM_RANGES-1:0][MAX_LENGTH*4-1:0] low;
    logic [NUM_RANGES-1:0][MAX_LENGTH*4-1:0] high;

    logic [SUM_SIZE-1:0] out;

    puzzle2 dut (
        .clk(clk),
        .rst_n(rst_n),
        .vld(vld),
        .low(low),
        .high(high),
        .out(out)
    );

    // Clock generation
    initial clk = 0;
    always #5 clk = ~clk;

    initial begin
		#20
        rst_n = 0;
        vld   = 0;
        for (int i = 0; i < NUM_RANGES; i++) begin
			low[i]  = 40'b0;
			high[i] = 40'b0;
		end
		
		
		#20
        rst_n = 1;
		
		
		#200

        // Load BCD low/high values

        low[0]  = 40'b0000000000000000000000000100010010000111;
        low[1]  = 40'b0000011101010101011101000101001000000111;
        low[2]  = 40'b0000100101010100100010010101100001001000;
        low[3]  = 40'b0000000000000100001101011000100000110010;
        low[4]  = 40'b0000000000000000000000000000000000010101;
        low[5]  = 40'b0000000000000000000000000000000000000001;
        low[6]  = 40'b0000000000001001000110011000100000001000;
        low[7]  = 40'b0000000000000000011001010111100110000001;
        low[8]  = 40'b0110001001010110000010011000001101000110;
        low[9]  = 40'b0000000000000000000000000000000101000010;
        low[10]  = 40'b0000000000010011000010010010010100101001;
        low[11]  = 40'b0000000010010110001000000001001010010110;
        low[12]  = 40'b0000000000011001011101100111001101000000;
        low[13]  = 40'b0000000000000010100000001001000000110110;
        low[14]  = 40'b0000000000000000001100110101100001010000;
        low[15]  = 40'b0000000000000000000101110010010000110111;
        low[16]  = 40'b0000000000000000011101100100010000110100;
        low[17]  = 40'b0000000000000000100100010000010101000011;
        low[18]  = 40'b0000000000000010000101000010000101111001;
        low[19]  = 40'b0000000000000110011001001001010101000101;
        low[20]  = 40'b0110010001100100010110000111100001001001;
        low[21]  = 40'b0000000000000000100001011000001110011001;
        low[22]  = 40'b0000000000000000000000000001001100101000;
        low[23]  = 40'b0000000000000000000001110010011110011000;
        low[24]  = 40'b0000000010001001011101110111011100011001;
        low[25]  = 40'b0000000010010001100010010001011110010010;
        low[26]  = 40'b0000000000000000000000000000001100010100;
        low[27]  = 40'b0000000000000000000000000000000001001000;
        low[28]  = 40'b0000000000000000010100100111100100000011;
        low[29]  = 40'b0000000000000000000000100100001001000000;

        high[0] = 40'b0000000000000000000000001001010110000001;
        high[1] = 40'b0000011101010101011101100110000010011001;
        high[2] = 40'b0000100101010101000001100011000100100100;
        high[3] = 40'b0000000000000100010010010111001100010101;
        high[4] = 40'b0000000000000000000000000000000001000111;
        high[5] = 40'b0000000000000000000000000000000000010010;
        high[6] = 40'b0000000000001001001001011000011101110001;
        high[7] = 40'b0000000000000000011101100010001001110101;
        high[8] = 40'b0110001001010110001100000011100001110010;
        high[9] = 40'b0000000000000000000000000000001010000010;
        high[10] = 40'b0000000000010011000101111001010100101000;
        high[11] = 40'b0000000010010110001101000001100001111001;
        high[12] = 40'b0000000000011001100100010110001101111000;
        high[13] = 40'b0000000000000010100000110000100001100010;
        high[14] = 40'b0000000000000000010010011001100110000110;
        high[15] = 40'b0000000000000000001100010101000101000100;
        high[16] = 40'b0000000000000000011110010011000100110011;
        high[17] = 40'b0000000000000001000010000010011001110000;
        high[18] = 40'b0000000000000010001001111001001000000011;
        high[19] = 40'b0000000000000110011100010011000010011000;
        high[20] = 40'b0110010001100100011001110111000000100100;
        high[21] = 40'b0000000000000000100100000100010010010001;
        high[22] = 40'b0000000000000000000000000100000000100001;
        high[23] = 40'b0000000000000000000101011001001000000110;
        high[24] = 40'b0000000010010000000000000101100000010010;
        high[25] = 40'b0000000010010001100100111000001001111001;
        high[26] = 40'b0000000000000000000000000000100101100011;
        high[27] = 40'b0000000000000000000000000000000100110000;
        high[28] = 40'b0000000000000000010110010100001101110000;
        high[29] = 40'b0000000000000000000001100000001000010010;


		#200
        vld   = 1;

        // Run long enough for DUT to complete internal accumulation
        #5000000;

        $display("\nDUT OUT = %0d (decimal)", out);
        $display("DUT OUT (hex) = %h", out);
        $display("DUT OUT (binary) = %b", out);

        $finish;
    end
	
	
initial begin
	/*
    $monitor(
        "T=%0t | clk=%0b rst_n=%0b vld=%0b | out=%0d low=%0d high=%0d num_q=%0d num_d=%0d num_vld_digit=%0d invalid=%0d sum_q=%0d sum_d=%0d done_q=%0d done_d=%0d cnt_q=%0d cnt_d=%0d direct_sum=%0d correct_sum=%0d num_to_binary=%0d all_range_sum_q=%0d",
        $time,
        clk, rst_n, vld,
        out,
        low[0],
        high[0],
        dut.num_q[0],
        dut.num_d[0],
		dut.num_vld_digit[0],
		dut.invalid_id[0],
        dut.sum_q[0],
        dut.sum_d[0],
        dut.done_q,
        dut.done_d,
        dut.cnt_q, dut.cnt_d,
        dut.direct_sum[0],
        dut.correct_sum[0],
        dut.num_to_binary[0],
        dut.all_range_sum_q,
        dut.all_range_sum_d
    );
	*/
	
	
	$monitor(
        "T=%0t | out=%0d low=%0d high=%0d num_q=%0d num_d=%0d num_vld_digit=%0d invalid=%0d sum_q=%0d sum_d=%0d done_q=%0d done_d=%0d cnt_q=%0d cnt_d=%0d direct_sum=%0d correct_sum=%0d num_to_binary=%0d all_range_sum_q=%0d",
        $time,
        out,
        low[0],
        high[0],
        dut.num_q[0],
        dut.num_d[0],
		dut.num_vld_digit[0],
		dut.invalid_id[0],
        dut.sum_q[0],
        dut.sum_d[0],
        dut.done_q,
        dut.done_d,
        dut.cnt_q, dut.cnt_d,
        dut.direct_sum[0],
        dut.correct_sum[0],
        dut.num_to_binary[0],
        dut.all_range_sum_q
    );
	

end

final begin
	// Print all 200 banks
	for (int i = 0; i < 30; i++) begin
		$display("sum[%0d] : %0d",
				i,
				dut.sum_q[i]
		);
	end
end


endmodule
